library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all; 
library std;    
use std.textio.all;
library work;
use work.pack_mips.all;
use work.txt_util.all;
library modelsim_lib;
use modelsim_lib.util.all;

entity sim_minimips is
end;

architecture bench of sim_minimips is

  component minimips is 
  port (
      clock    : in std_logic;
      reset    : in std_logic;
      ram_req  : out std_logic;
      ram_adr  : out bus32;
      ram_r_w  : out std_logic;
      ram_data : inout bus32;
      ram_ack  : in std_logic;
      -- Caco
      --mem_data_in  : in bus32;
      mem_data_out : out bus32;
      --
      it_mat   : in std_logic
  );
  end component;
  

  component ram is
    generic (mem_size : natural := 8192;
             latency : time := 10 ns);
    port(
        req        	: in std_logic;
        adr        	: in bus32;
        -- Caco
        mem_data_in  : in bus32;
--        mem_data_out : out bus32;
        --
        data_inout 	: inout bus32;
        r_w        	: in std_logic;
        ready      	: out std_logic;
		reset		: in std_logic;
		clock		: in std_logic
	);

  end component;


  signal clock : std_logic;
  signal reset : std_logic;
  signal it_mat : std_logic := '0';
  -- Connexion with the Ram
  signal ram_req : std_logic;
  signal ram_adr : bus32;
  signal ram_r_w : std_logic;
  signal ram_data : bus32;
  signal ram_data_temp : bus32;
  signal ram_rdy : std_logic;
  signal mem_data_out_in : bus32;
  signal end_of_execution : std_logic := '0';
  signal debug1 : std_logic := '0'; 
  
  signal clock_g : std_logic;
  signal reset_g : std_logic;
  signal it_mat_g : std_logic := '0';
  -- Connexion with the Ram
  signal ram_req_g : std_logic;
  signal ram_adr_g : bus32;
  signal ram_r_w_g : std_logic;
  signal ram_data_g : bus32;
  signal ram_data_temp_g : bus32;
  signal ram_rdy_g : std_logic;
  signal mem_data_out_in_g : bus32;
  signal end_of_execution_g : std_logic := '0';
  signal debug1_g : std_logic := '0'; 
  
  
 signal control_uut : std_logic_vector (1 to 911); -- tamanho igual a lista de sinais
 signal control_gold : std_logic_vector (1 to 911); -- tamanho igual a lista de sinais

	type list_string1 is array (natural range <> ) of string(1 to 59);
   constant control_signals_uut : list_string1(1 to 911) := 
(
"/sim_minimips/u_minimips/u1_pf/suivant(0)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(1)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(2)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(3)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(4)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(5)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(6)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(7)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(8)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(9)                  ",
"/sim_minimips/u_minimips/u1_pf/suivant(10)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(11)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(12)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(13)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(14)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(15)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(16)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(17)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(18)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(19)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(20)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(21)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(22)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(23)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(24)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(25)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(26)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(27)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(28)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(29)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(30)                 ",
"/sim_minimips/u_minimips/u1_pf/suivant(31)                 ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(0)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(1)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(2)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(3)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(4)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(5)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(6)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(7)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(8)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(9)               ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(10)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(11)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(12)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(13)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(14)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(15)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(16)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(17)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(18)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(19)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(20)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(21)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(22)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(23)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(24)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(25)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(26)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(27)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(28)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(29)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(30)              ",
"/sim_minimips/u_minimips/u1_pf/pc_interne(31)              ",
"/sim_minimips/u_minimips/u1_pf/lock                        ",
"/sim_minimips/u_minimips/clock                             ",
"/sim_minimips/u_minimips/reset                             ",
"/sim_minimips/u_minimips/ram_req                           ",
"/sim_minimips/u_minimips/ram_adr(0)                        ",
"/sim_minimips/u_minimips/ram_adr(1)                        ",
"/sim_minimips/u_minimips/ram_adr(2)                        ",
"/sim_minimips/u_minimips/ram_adr(3)                        ",
"/sim_minimips/u_minimips/ram_adr(4)                        ",
"/sim_minimips/u_minimips/ram_adr(5)                        ",
"/sim_minimips/u_minimips/ram_adr(6)                        ",
"/sim_minimips/u_minimips/ram_adr(7)                        ",
"/sim_minimips/u_minimips/ram_adr(8)                        ",
"/sim_minimips/u_minimips/ram_adr(9)                        ",
"/sim_minimips/u_minimips/ram_adr(10)                       ",
"/sim_minimips/u_minimips/ram_adr(11)                       ",
"/sim_minimips/u_minimips/ram_adr(12)                       ",
"/sim_minimips/u_minimips/ram_adr(13)                       ",
"/sim_minimips/u_minimips/ram_adr(14)                       ",
"/sim_minimips/u_minimips/ram_adr(15)                       ",
"/sim_minimips/u_minimips/ram_adr(16)                       ",
"/sim_minimips/u_minimips/ram_adr(17)                       ",
"/sim_minimips/u_minimips/ram_adr(18)                       ",
"/sim_minimips/u_minimips/ram_adr(19)                       ",
"/sim_minimips/u_minimips/ram_adr(20)                       ",
"/sim_minimips/u_minimips/ram_adr(21)                       ",
"/sim_minimips/u_minimips/ram_adr(22)                       ",
"/sim_minimips/u_minimips/ram_adr(23)                       ",
"/sim_minimips/u_minimips/ram_adr(24)                       ",
"/sim_minimips/u_minimips/ram_adr(25)                       ",
"/sim_minimips/u_minimips/ram_adr(26)                       ",
"/sim_minimips/u_minimips/ram_adr(27)                       ",
"/sim_minimips/u_minimips/ram_adr(28)                       ",
"/sim_minimips/u_minimips/ram_adr(29)                       ",
"/sim_minimips/u_minimips/ram_adr(30)                       ",
"/sim_minimips/u_minimips/ram_adr(31)                       ",
"/sim_minimips/u_minimips/ram_r_w                           ",
"/sim_minimips/u_minimips/ram_ack                           ",
"/sim_minimips/u_minimips/it_mat                            ",
"/sim_minimips/u_minimips/stop_all                          ",
"/sim_minimips/u_minimips/it_mat_clk                        ",
"/sim_minimips/u_minimips/pf_pc(0)                          ",
"/sim_minimips/u_minimips/pf_pc(1)                          ",
"/sim_minimips/u_minimips/pf_pc(2)                          ",
"/sim_minimips/u_minimips/pf_pc(3)                          ",
"/sim_minimips/u_minimips/pf_pc(4)                          ",
"/sim_minimips/u_minimips/pf_pc(5)                          ",
"/sim_minimips/u_minimips/pf_pc(6)                          ",
"/sim_minimips/u_minimips/pf_pc(7)                          ",
"/sim_minimips/u_minimips/pf_pc(8)                          ",
"/sim_minimips/u_minimips/pf_pc(9)                          ",
"/sim_minimips/u_minimips/pf_pc(10)                         ",
"/sim_minimips/u_minimips/pf_pc(11)                         ",
"/sim_minimips/u_minimips/pf_pc(12)                         ",
"/sim_minimips/u_minimips/pf_pc(13)                         ",
"/sim_minimips/u_minimips/pf_pc(14)                         ",
"/sim_minimips/u_minimips/pf_pc(15)                         ",
"/sim_minimips/u_minimips/pf_pc(16)                         ",
"/sim_minimips/u_minimips/pf_pc(17)                         ",
"/sim_minimips/u_minimips/pf_pc(18)                         ",
"/sim_minimips/u_minimips/pf_pc(19)                         ",
"/sim_minimips/u_minimips/pf_pc(20)                         ",
"/sim_minimips/u_minimips/pf_pc(21)                         ",
"/sim_minimips/u_minimips/pf_pc(22)                         ",
"/sim_minimips/u_minimips/pf_pc(23)                         ",
"/sim_minimips/u_minimips/pf_pc(24)                         ",
"/sim_minimips/u_minimips/pf_pc(25)                         ",
"/sim_minimips/u_minimips/pf_pc(26)                         ",
"/sim_minimips/u_minimips/pf_pc(27)                         ",
"/sim_minimips/u_minimips/pf_pc(28)                         ",
"/sim_minimips/u_minimips/pf_pc(29)                         ",
"/sim_minimips/u_minimips/pf_pc(30)                         ",
"/sim_minimips/u_minimips/pf_pc(31)                         ",
"/sim_minimips/u_minimips/cte_instr(0)                      ",
"/sim_minimips/u_minimips/cte_instr(1)                      ",
"/sim_minimips/u_minimips/cte_instr(2)                      ",
"/sim_minimips/u_minimips/cte_instr(3)                      ",
"/sim_minimips/u_minimips/cte_instr(4)                      ",
"/sim_minimips/u_minimips/cte_instr(5)                      ",
"/sim_minimips/u_minimips/cte_instr(6)                      ",
"/sim_minimips/u_minimips/cte_instr(7)                      ",
"/sim_minimips/u_minimips/cte_instr(8)                      ",
"/sim_minimips/u_minimips/cte_instr(9)                      ",
"/sim_minimips/u_minimips/cte_instr(10)                     ",
"/sim_minimips/u_minimips/cte_instr(11)                     ",
"/sim_minimips/u_minimips/cte_instr(12)                     ",
"/sim_minimips/u_minimips/cte_instr(13)                     ",
"/sim_minimips/u_minimips/cte_instr(14)                     ",
"/sim_minimips/u_minimips/cte_instr(15)                     ",
"/sim_minimips/u_minimips/cte_instr(16)                     ",
"/sim_minimips/u_minimips/cte_instr(17)                     ",
"/sim_minimips/u_minimips/cte_instr(18)                     ",
"/sim_minimips/u_minimips/cte_instr(19)                     ",
"/sim_minimips/u_minimips/cte_instr(20)                     ",
"/sim_minimips/u_minimips/cte_instr(21)                     ",
"/sim_minimips/u_minimips/cte_instr(22)                     ",
"/sim_minimips/u_minimips/cte_instr(23)                     ",
"/sim_minimips/u_minimips/cte_instr(24)                     ",
"/sim_minimips/u_minimips/cte_instr(25)                     ",
"/sim_minimips/u_minimips/cte_instr(26)                     ",
"/sim_minimips/u_minimips/cte_instr(27)                     ",
"/sim_minimips/u_minimips/cte_instr(28)                     ",
"/sim_minimips/u_minimips/cte_instr(29)                     ",
"/sim_minimips/u_minimips/cte_instr(30)                     ",
"/sim_minimips/u_minimips/cte_instr(31)                     ",
"/sim_minimips/u_minimips/etc_adr(0)                        ",
"/sim_minimips/u_minimips/etc_adr(1)                        ",
"/sim_minimips/u_minimips/etc_adr(2)                        ",
"/sim_minimips/u_minimips/etc_adr(3)                        ",
"/sim_minimips/u_minimips/etc_adr(4)                        ",
"/sim_minimips/u_minimips/etc_adr(5)                        ",
"/sim_minimips/u_minimips/etc_adr(6)                        ",
"/sim_minimips/u_minimips/etc_adr(7)                        ",
"/sim_minimips/u_minimips/etc_adr(8)                        ",
"/sim_minimips/u_minimips/etc_adr(9)                        ",
"/sim_minimips/u_minimips/etc_adr(10)                       ",
"/sim_minimips/u_minimips/etc_adr(11)                       ",
"/sim_minimips/u_minimips/etc_adr(12)                       ",
"/sim_minimips/u_minimips/etc_adr(13)                       ",
"/sim_minimips/u_minimips/etc_adr(14)                       ",
"/sim_minimips/u_minimips/etc_adr(15)                       ",
"/sim_minimips/u_minimips/etc_adr(16)                       ",
"/sim_minimips/u_minimips/etc_adr(17)                       ",
"/sim_minimips/u_minimips/etc_adr(18)                       ",
"/sim_minimips/u_minimips/etc_adr(19)                       ",
"/sim_minimips/u_minimips/etc_adr(20)                       ",
"/sim_minimips/u_minimips/etc_adr(21)                       ",
"/sim_minimips/u_minimips/etc_adr(22)                       ",
"/sim_minimips/u_minimips/etc_adr(23)                       ",
"/sim_minimips/u_minimips/etc_adr(24)                       ",
"/sim_minimips/u_minimips/etc_adr(25)                       ",
"/sim_minimips/u_minimips/etc_adr(26)                       ",
"/sim_minimips/u_minimips/etc_adr(27)                       ",
"/sim_minimips/u_minimips/etc_adr(28)                       ",
"/sim_minimips/u_minimips/etc_adr(29)                       ",
"/sim_minimips/u_minimips/etc_adr(30)                       ",
"/sim_minimips/u_minimips/etc_adr(31)                       ",
"/sim_minimips/u_minimips/ei_instr(0)                       ",
"/sim_minimips/u_minimips/ei_instr(1)                       ",
"/sim_minimips/u_minimips/ei_instr(2)                       ",
"/sim_minimips/u_minimips/ei_instr(3)                       ",
"/sim_minimips/u_minimips/ei_instr(4)                       ",
"/sim_minimips/u_minimips/ei_instr(5)                       ",
"/sim_minimips/u_minimips/ei_instr(6)                       ",
"/sim_minimips/u_minimips/ei_instr(7)                       ",
"/sim_minimips/u_minimips/ei_instr(8)                       ",
"/sim_minimips/u_minimips/ei_instr(9)                       ",
"/sim_minimips/u_minimips/ei_instr(10)                      ",
"/sim_minimips/u_minimips/ei_instr(11)                      ",
"/sim_minimips/u_minimips/ei_instr(12)                      ",
"/sim_minimips/u_minimips/ei_instr(13)                      ",
"/sim_minimips/u_minimips/ei_instr(14)                      ",
"/sim_minimips/u_minimips/ei_instr(15)                      ",
"/sim_minimips/u_minimips/ei_instr(16)                      ",
"/sim_minimips/u_minimips/ei_instr(17)                      ",
"/sim_minimips/u_minimips/ei_instr(18)                      ",
"/sim_minimips/u_minimips/ei_instr(19)                      ",
"/sim_minimips/u_minimips/ei_instr(20)                      ",
"/sim_minimips/u_minimips/ei_instr(21)                      ",
"/sim_minimips/u_minimips/ei_instr(22)                      ",
"/sim_minimips/u_minimips/ei_instr(23)                      ",
"/sim_minimips/u_minimips/ei_instr(24)                      ",
"/sim_minimips/u_minimips/ei_instr(25)                      ",
"/sim_minimips/u_minimips/ei_instr(26)                      ",
"/sim_minimips/u_minimips/ei_instr(27)                      ",
"/sim_minimips/u_minimips/ei_instr(28)                      ",
"/sim_minimips/u_minimips/ei_instr(29)                      ",
"/sim_minimips/u_minimips/ei_instr(30)                      ",
"/sim_minimips/u_minimips/ei_instr(31)                      ",
"/sim_minimips/u_minimips/ei_adr(0)                         ",
"/sim_minimips/u_minimips/ei_adr(1)                         ",
"/sim_minimips/u_minimips/ei_adr(2)                         ",
"/sim_minimips/u_minimips/ei_adr(3)                         ",
"/sim_minimips/u_minimips/ei_adr(4)                         ",
"/sim_minimips/u_minimips/ei_adr(5)                         ",
"/sim_minimips/u_minimips/ei_adr(6)                         ",
"/sim_minimips/u_minimips/ei_adr(7)                         ",
"/sim_minimips/u_minimips/ei_adr(8)                         ",
"/sim_minimips/u_minimips/ei_adr(9)                         ",
"/sim_minimips/u_minimips/ei_adr(10)                        ",
"/sim_minimips/u_minimips/ei_adr(11)                        ",
"/sim_minimips/u_minimips/ei_adr(12)                        ",
"/sim_minimips/u_minimips/ei_adr(13)                        ",
"/sim_minimips/u_minimips/ei_adr(14)                        ",
"/sim_minimips/u_minimips/ei_adr(15)                        ",
"/sim_minimips/u_minimips/ei_adr(16)                        ",
"/sim_minimips/u_minimips/ei_adr(17)                        ",
"/sim_minimips/u_minimips/ei_adr(18)                        ",
"/sim_minimips/u_minimips/ei_adr(19)                        ",
"/sim_minimips/u_minimips/ei_adr(20)                        ",
"/sim_minimips/u_minimips/ei_adr(21)                        ",
"/sim_minimips/u_minimips/ei_adr(22)                        ",
"/sim_minimips/u_minimips/ei_adr(23)                        ",
"/sim_minimips/u_minimips/ei_adr(24)                        ",
"/sim_minimips/u_minimips/ei_adr(25)                        ",
"/sim_minimips/u_minimips/ei_adr(26)                        ",
"/sim_minimips/u_minimips/ei_adr(27)                        ",
"/sim_minimips/u_minimips/ei_adr(28)                        ",
"/sim_minimips/u_minimips/ei_adr(29)                        ",
"/sim_minimips/u_minimips/ei_adr(30)                        ",
"/sim_minimips/u_minimips/ei_adr(31)                        ",
"/sim_minimips/u_minimips/ei_it_ok                          ",
"/sim_minimips/u_minimips/adr_reg1(0)                       ",
"/sim_minimips/u_minimips/adr_reg1(1)                       ",
"/sim_minimips/u_minimips/adr_reg1(2)                       ",
"/sim_minimips/u_minimips/adr_reg1(3)                       ",
"/sim_minimips/u_minimips/adr_reg1(4)                       ",
"/sim_minimips/u_minimips/adr_reg1(5)                       ",
"/sim_minimips/u_minimips/adr_reg2(0)                       ",
"/sim_minimips/u_minimips/adr_reg2(1)                       ",
"/sim_minimips/u_minimips/adr_reg2(2)                       ",
"/sim_minimips/u_minimips/adr_reg2(3)                       ",
"/sim_minimips/u_minimips/adr_reg2(4)                       ",
"/sim_minimips/u_minimips/adr_reg2(5)                       ",
"/sim_minimips/u_minimips/use1                              ",
"/sim_minimips/u_minimips/use2                              ",
"/sim_minimips/u_minimips/alea                              ",
"/sim_minimips/u_minimips/di_bra                            ",
"/sim_minimips/u_minimips/di_link                           ",
"/sim_minimips/u_minimips/di_code_ual(0)                    ",
"/sim_minimips/u_minimips/di_code_ual(1)                    ",
"/sim_minimips/u_minimips/di_code_ual(2)                    ",
"/sim_minimips/u_minimips/di_code_ual(3)                    ",
"/sim_minimips/u_minimips/di_code_ual(4)                    ",
"/sim_minimips/u_minimips/di_code_ual(5)                    ",
"/sim_minimips/u_minimips/di_code_ual(6)                    ",
"/sim_minimips/u_minimips/di_code_ual(7)                    ",
"/sim_minimips/u_minimips/di_code_ual(8)                    ",
"/sim_minimips/u_minimips/di_code_ual(9)                    ",
"/sim_minimips/u_minimips/di_code_ual(10)                   ",
"/sim_minimips/u_minimips/di_code_ual(11)                   ",
"/sim_minimips/u_minimips/di_code_ual(12)                   ",
"/sim_minimips/u_minimips/di_code_ual(13)                   ",
"/sim_minimips/u_minimips/di_code_ual(14)                   ",
"/sim_minimips/u_minimips/di_code_ual(15)                   ",
"/sim_minimips/u_minimips/di_code_ual(16)                   ",
"/sim_minimips/u_minimips/di_code_ual(17)                   ",
"/sim_minimips/u_minimips/di_code_ual(18)                   ",
"/sim_minimips/u_minimips/di_code_ual(19)                   ",
"/sim_minimips/u_minimips/di_code_ual(20)                   ",
"/sim_minimips/u_minimips/di_code_ual(21)                   ",
"/sim_minimips/u_minimips/di_code_ual(22)                   ",
"/sim_minimips/u_minimips/di_code_ual(23)                   ",
"/sim_minimips/u_minimips/di_code_ual(24)                   ",
"/sim_minimips/u_minimips/di_code_ual(25)                   ",
"/sim_minimips/u_minimips/di_code_ual(26)                   ",
"/sim_minimips/u_minimips/di_code_ual(27)                   ",
"/sim_minimips/u_minimips/di_offset(0)                      ",
"/sim_minimips/u_minimips/di_offset(1)                      ",
"/sim_minimips/u_minimips/di_offset(2)                      ",
"/sim_minimips/u_minimips/di_offset(3)                      ",
"/sim_minimips/u_minimips/di_offset(4)                      ",
"/sim_minimips/u_minimips/di_offset(5)                      ",
"/sim_minimips/u_minimips/di_offset(6)                      ",
"/sim_minimips/u_minimips/di_offset(7)                      ",
"/sim_minimips/u_minimips/di_offset(8)                      ",
"/sim_minimips/u_minimips/di_offset(9)                      ",
"/sim_minimips/u_minimips/di_offset(10)                     ",
"/sim_minimips/u_minimips/di_offset(11)                     ",
"/sim_minimips/u_minimips/di_offset(12)                     ",
"/sim_minimips/u_minimips/di_offset(13)                     ",
"/sim_minimips/u_minimips/di_offset(14)                     ",
"/sim_minimips/u_minimips/di_offset(15)                     ",
"/sim_minimips/u_minimips/di_offset(16)                     ",
"/sim_minimips/u_minimips/di_offset(17)                     ",
"/sim_minimips/u_minimips/di_offset(18)                     ",
"/sim_minimips/u_minimips/di_offset(19)                     ",
"/sim_minimips/u_minimips/di_offset(20)                     ",
"/sim_minimips/u_minimips/di_offset(21)                     ",
"/sim_minimips/u_minimips/di_offset(22)                     ",
"/sim_minimips/u_minimips/di_offset(23)                     ",
"/sim_minimips/u_minimips/di_offset(24)                     ",
"/sim_minimips/u_minimips/di_offset(25)                     ",
"/sim_minimips/u_minimips/di_offset(26)                     ",
"/sim_minimips/u_minimips/di_offset(27)                     ",
"/sim_minimips/u_minimips/di_offset(28)                     ",
"/sim_minimips/u_minimips/di_offset(29)                     ",
"/sim_minimips/u_minimips/di_offset(30)                     ",
"/sim_minimips/u_minimips/di_offset(31)                     ",
"/sim_minimips/u_minimips/di_adr_reg_dest(0)                ",
"/sim_minimips/u_minimips/di_adr_reg_dest(1)                ",
"/sim_minimips/u_minimips/di_adr_reg_dest(2)                ",
"/sim_minimips/u_minimips/di_adr_reg_dest(3)                ",
"/sim_minimips/u_minimips/di_adr_reg_dest(4)                ",
"/sim_minimips/u_minimips/di_adr_reg_dest(5)                ",
"/sim_minimips/u_minimips/di_ecr_reg                        ",
"/sim_minimips/u_minimips/di_mode                           ",
"/sim_minimips/u_minimips/di_op_mem                         ",
"/sim_minimips/u_minimips/di_r_w                            ",
"/sim_minimips/u_minimips/di_adr(0)                         ",
"/sim_minimips/u_minimips/di_adr(1)                         ",
"/sim_minimips/u_minimips/di_adr(2)                         ",
"/sim_minimips/u_minimips/di_adr(3)                         ",
"/sim_minimips/u_minimips/di_adr(4)                         ",
"/sim_minimips/u_minimips/di_adr(5)                         ",
"/sim_minimips/u_minimips/di_adr(6)                         ",
"/sim_minimips/u_minimips/di_adr(7)                         ",
"/sim_minimips/u_minimips/di_adr(8)                         ",
"/sim_minimips/u_minimips/di_adr(9)                         ",
"/sim_minimips/u_minimips/di_adr(10)                        ",
"/sim_minimips/u_minimips/di_adr(11)                        ",
"/sim_minimips/u_minimips/di_adr(12)                        ",
"/sim_minimips/u_minimips/di_adr(13)                        ",
"/sim_minimips/u_minimips/di_adr(14)                        ",
"/sim_minimips/u_minimips/di_adr(15)                        ",
"/sim_minimips/u_minimips/di_adr(16)                        ",
"/sim_minimips/u_minimips/di_adr(17)                        ",
"/sim_minimips/u_minimips/di_adr(18)                        ",
"/sim_minimips/u_minimips/di_adr(19)                        ",
"/sim_minimips/u_minimips/di_adr(20)                        ",
"/sim_minimips/u_minimips/di_adr(21)                        ",
"/sim_minimips/u_minimips/di_adr(22)                        ",
"/sim_minimips/u_minimips/di_adr(23)                        ",
"/sim_minimips/u_minimips/di_adr(24)                        ",
"/sim_minimips/u_minimips/di_adr(25)                        ",
"/sim_minimips/u_minimips/di_adr(26)                        ",
"/sim_minimips/u_minimips/di_adr(27)                        ",
"/sim_minimips/u_minimips/di_adr(28)                        ",
"/sim_minimips/u_minimips/di_adr(29)                        ",
"/sim_minimips/u_minimips/di_adr(30)                        ",
"/sim_minimips/u_minimips/di_adr(31)                        ",
"/sim_minimips/u_minimips/di_exc_cause(0)                   ",
"/sim_minimips/u_minimips/di_exc_cause(1)                   ",
"/sim_minimips/u_minimips/di_exc_cause(2)                   ",
"/sim_minimips/u_minimips/di_exc_cause(3)                   ",
"/sim_minimips/u_minimips/di_exc_cause(4)                   ",
"/sim_minimips/u_minimips/di_exc_cause(5)                   ",
"/sim_minimips/u_minimips/di_exc_cause(6)                   ",
"/sim_minimips/u_minimips/di_exc_cause(7)                   ",
"/sim_minimips/u_minimips/di_exc_cause(8)                   ",
"/sim_minimips/u_minimips/di_exc_cause(9)                   ",
"/sim_minimips/u_minimips/di_exc_cause(10)                  ",
"/sim_minimips/u_minimips/di_exc_cause(11)                  ",
"/sim_minimips/u_minimips/di_exc_cause(12)                  ",
"/sim_minimips/u_minimips/di_exc_cause(13)                  ",
"/sim_minimips/u_minimips/di_exc_cause(14)                  ",
"/sim_minimips/u_minimips/di_exc_cause(15)                  ",
"/sim_minimips/u_minimips/di_exc_cause(16)                  ",
"/sim_minimips/u_minimips/di_exc_cause(17)                  ",
"/sim_minimips/u_minimips/di_exc_cause(18)                  ",
"/sim_minimips/u_minimips/di_exc_cause(19)                  ",
"/sim_minimips/u_minimips/di_exc_cause(20)                  ",
"/sim_minimips/u_minimips/di_exc_cause(21)                  ",
"/sim_minimips/u_minimips/di_exc_cause(22)                  ",
"/sim_minimips/u_minimips/di_exc_cause(23)                  ",
"/sim_minimips/u_minimips/di_exc_cause(24)                  ",
"/sim_minimips/u_minimips/di_exc_cause(25)                  ",
"/sim_minimips/u_minimips/di_exc_cause(26)                  ",
"/sim_minimips/u_minimips/di_exc_cause(27)                  ",
"/sim_minimips/u_minimips/di_exc_cause(28)                  ",
"/sim_minimips/u_minimips/di_exc_cause(29)                  ",
"/sim_minimips/u_minimips/di_exc_cause(30)                  ",
"/sim_minimips/u_minimips/di_exc_cause(31)                  ",
"/sim_minimips/u_minimips/di_level(0)                       ",
"/sim_minimips/u_minimips/di_level(1)                       ",
"/sim_minimips/u_minimips/di_it_ok                          ",
"/sim_minimips/u_minimips/ex_adr(0)                         ",
"/sim_minimips/u_minimips/ex_adr(1)                         ",
"/sim_minimips/u_minimips/ex_adr(2)                         ",
"/sim_minimips/u_minimips/ex_adr(3)                         ",
"/sim_minimips/u_minimips/ex_adr(4)                         ",
"/sim_minimips/u_minimips/ex_adr(5)                         ",
"/sim_minimips/u_minimips/ex_adr(6)                         ",
"/sim_minimips/u_minimips/ex_adr(7)                         ",
"/sim_minimips/u_minimips/ex_adr(8)                         ",
"/sim_minimips/u_minimips/ex_adr(9)                         ",
"/sim_minimips/u_minimips/ex_adr(10)                        ",
"/sim_minimips/u_minimips/ex_adr(11)                        ",
"/sim_minimips/u_minimips/ex_adr(12)                        ",
"/sim_minimips/u_minimips/ex_adr(13)                        ",
"/sim_minimips/u_minimips/ex_adr(14)                        ",
"/sim_minimips/u_minimips/ex_adr(15)                        ",
"/sim_minimips/u_minimips/ex_adr(16)                        ",
"/sim_minimips/u_minimips/ex_adr(17)                        ",
"/sim_minimips/u_minimips/ex_adr(18)                        ",
"/sim_minimips/u_minimips/ex_adr(19)                        ",
"/sim_minimips/u_minimips/ex_adr(20)                        ",
"/sim_minimips/u_minimips/ex_adr(21)                        ",
"/sim_minimips/u_minimips/ex_adr(22)                        ",
"/sim_minimips/u_minimips/ex_adr(23)                        ",
"/sim_minimips/u_minimips/ex_adr(24)                        ",
"/sim_minimips/u_minimips/ex_adr(25)                        ",
"/sim_minimips/u_minimips/ex_adr(26)                        ",
"/sim_minimips/u_minimips/ex_adr(27)                        ",
"/sim_minimips/u_minimips/ex_adr(28)                        ",
"/sim_minimips/u_minimips/ex_adr(29)                        ",
"/sim_minimips/u_minimips/ex_adr(30)                        ",
"/sim_minimips/u_minimips/ex_adr(31)                        ",
"/sim_minimips/u_minimips/ex_bra_confirm                    ",
"/sim_minimips/u_minimips/ex_adresse(0)                     ",
"/sim_minimips/u_minimips/ex_adresse(1)                     ",
"/sim_minimips/u_minimips/ex_adresse(2)                     ",
"/sim_minimips/u_minimips/ex_adresse(3)                     ",
"/sim_minimips/u_minimips/ex_adresse(4)                     ",
"/sim_minimips/u_minimips/ex_adresse(5)                     ",
"/sim_minimips/u_minimips/ex_adresse(6)                     ",
"/sim_minimips/u_minimips/ex_adresse(7)                     ",
"/sim_minimips/u_minimips/ex_adresse(8)                     ",
"/sim_minimips/u_minimips/ex_adresse(9)                     ",
"/sim_minimips/u_minimips/ex_adresse(10)                    ",
"/sim_minimips/u_minimips/ex_adresse(11)                    ",
"/sim_minimips/u_minimips/ex_adresse(12)                    ",
"/sim_minimips/u_minimips/ex_adresse(13)                    ",
"/sim_minimips/u_minimips/ex_adresse(14)                    ",
"/sim_minimips/u_minimips/ex_adresse(15)                    ",
"/sim_minimips/u_minimips/ex_adresse(16)                    ",
"/sim_minimips/u_minimips/ex_adresse(17)                    ",
"/sim_minimips/u_minimips/ex_adresse(18)                    ",
"/sim_minimips/u_minimips/ex_adresse(19)                    ",
"/sim_minimips/u_minimips/ex_adresse(20)                    ",
"/sim_minimips/u_minimips/ex_adresse(21)                    ",
"/sim_minimips/u_minimips/ex_adresse(22)                    ",
"/sim_minimips/u_minimips/ex_adresse(23)                    ",
"/sim_minimips/u_minimips/ex_adresse(24)                    ",
"/sim_minimips/u_minimips/ex_adresse(25)                    ",
"/sim_minimips/u_minimips/ex_adresse(26)                    ",
"/sim_minimips/u_minimips/ex_adresse(27)                    ",
"/sim_minimips/u_minimips/ex_adresse(28)                    ",
"/sim_minimips/u_minimips/ex_adresse(29)                    ",
"/sim_minimips/u_minimips/ex_adresse(30)                    ",
"/sim_minimips/u_minimips/ex_adresse(31)                    ",
"/sim_minimips/u_minimips/ex_adr_reg_dest(0)                ",
"/sim_minimips/u_minimips/ex_adr_reg_dest(1)                ",
"/sim_minimips/u_minimips/ex_adr_reg_dest(2)                ",
"/sim_minimips/u_minimips/ex_adr_reg_dest(3)                ",
"/sim_minimips/u_minimips/ex_adr_reg_dest(4)                ",
"/sim_minimips/u_minimips/ex_adr_reg_dest(5)                ",
"/sim_minimips/u_minimips/ex_ecr_reg                        ",
"/sim_minimips/u_minimips/ex_op_mem                         ",
"/sim_minimips/u_minimips/ex_r_w                            ",
"/sim_minimips/u_minimips/ex_exc_cause(0)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(1)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(2)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(3)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(4)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(5)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(6)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(7)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(8)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(9)                   ",
"/sim_minimips/u_minimips/ex_exc_cause(10)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(11)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(12)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(13)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(14)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(15)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(16)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(17)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(18)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(19)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(20)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(21)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(22)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(23)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(24)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(25)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(26)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(27)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(28)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(29)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(30)                  ",
"/sim_minimips/u_minimips/ex_exc_cause(31)                  ",
"/sim_minimips/u_minimips/ex_level(0)                       ",
"/sim_minimips/u_minimips/ex_level(1)                       ",
"/sim_minimips/u_minimips/ex_it_ok                          ",
"/sim_minimips/u_minimips/mtc_adr(0)                        ",
"/sim_minimips/u_minimips/mtc_adr(1)                        ",
"/sim_minimips/u_minimips/mtc_adr(2)                        ",
"/sim_minimips/u_minimips/mtc_adr(3)                        ",
"/sim_minimips/u_minimips/mtc_adr(4)                        ",
"/sim_minimips/u_minimips/mtc_adr(5)                        ",
"/sim_minimips/u_minimips/mtc_adr(6)                        ",
"/sim_minimips/u_minimips/mtc_adr(7)                        ",
"/sim_minimips/u_minimips/mtc_adr(8)                        ",
"/sim_minimips/u_minimips/mtc_adr(9)                        ",
"/sim_minimips/u_minimips/mtc_adr(10)                       ",
"/sim_minimips/u_minimips/mtc_adr(11)                       ",
"/sim_minimips/u_minimips/mtc_adr(12)                       ",
"/sim_minimips/u_minimips/mtc_adr(13)                       ",
"/sim_minimips/u_minimips/mtc_adr(14)                       ",
"/sim_minimips/u_minimips/mtc_adr(15)                       ",
"/sim_minimips/u_minimips/mtc_adr(16)                       ",
"/sim_minimips/u_minimips/mtc_adr(17)                       ",
"/sim_minimips/u_minimips/mtc_adr(18)                       ",
"/sim_minimips/u_minimips/mtc_adr(19)                       ",
"/sim_minimips/u_minimips/mtc_adr(20)                       ",
"/sim_minimips/u_minimips/mtc_adr(21)                       ",
"/sim_minimips/u_minimips/mtc_adr(22)                       ",
"/sim_minimips/u_minimips/mtc_adr(23)                       ",
"/sim_minimips/u_minimips/mtc_adr(24)                       ",
"/sim_minimips/u_minimips/mtc_adr(25)                       ",
"/sim_minimips/u_minimips/mtc_adr(26)                       ",
"/sim_minimips/u_minimips/mtc_adr(27)                       ",
"/sim_minimips/u_minimips/mtc_adr(28)                       ",
"/sim_minimips/u_minimips/mtc_adr(29)                       ",
"/sim_minimips/u_minimips/mtc_adr(30)                       ",
"/sim_minimips/u_minimips/mtc_adr(31)                       ",
"/sim_minimips/u_minimips/mtc_r_w                           ",
"/sim_minimips/u_minimips/mtc_req                           ",
"/sim_minimips/u_minimips/mem_adr(0)                        ",
"/sim_minimips/u_minimips/mem_adr(1)                        ",
"/sim_minimips/u_minimips/mem_adr(2)                        ",
"/sim_minimips/u_minimips/mem_adr(3)                        ",
"/sim_minimips/u_minimips/mem_adr(4)                        ",
"/sim_minimips/u_minimips/mem_adr(5)                        ",
"/sim_minimips/u_minimips/mem_adr(6)                        ",
"/sim_minimips/u_minimips/mem_adr(7)                        ",
"/sim_minimips/u_minimips/mem_adr(8)                        ",
"/sim_minimips/u_minimips/mem_adr(9)                        ",
"/sim_minimips/u_minimips/mem_adr(10)                       ",
"/sim_minimips/u_minimips/mem_adr(11)                       ",
"/sim_minimips/u_minimips/mem_adr(12)                       ",
"/sim_minimips/u_minimips/mem_adr(13)                       ",
"/sim_minimips/u_minimips/mem_adr(14)                       ",
"/sim_minimips/u_minimips/mem_adr(15)                       ",
"/sim_minimips/u_minimips/mem_adr(16)                       ",
"/sim_minimips/u_minimips/mem_adr(17)                       ",
"/sim_minimips/u_minimips/mem_adr(18)                       ",
"/sim_minimips/u_minimips/mem_adr(19)                       ",
"/sim_minimips/u_minimips/mem_adr(20)                       ",
"/sim_minimips/u_minimips/mem_adr(21)                       ",
"/sim_minimips/u_minimips/mem_adr(22)                       ",
"/sim_minimips/u_minimips/mem_adr(23)                       ",
"/sim_minimips/u_minimips/mem_adr(24)                       ",
"/sim_minimips/u_minimips/mem_adr(25)                       ",
"/sim_minimips/u_minimips/mem_adr(26)                       ",
"/sim_minimips/u_minimips/mem_adr(27)                       ",
"/sim_minimips/u_minimips/mem_adr(28)                       ",
"/sim_minimips/u_minimips/mem_adr(29)                       ",
"/sim_minimips/u_minimips/mem_adr(30)                       ",
"/sim_minimips/u_minimips/mem_adr(31)                       ",
"/sim_minimips/u_minimips/mem_adr_reg_dest(0)               ",
"/sim_minimips/u_minimips/mem_adr_reg_dest(1)               ",
"/sim_minimips/u_minimips/mem_adr_reg_dest(2)               ",
"/sim_minimips/u_minimips/mem_adr_reg_dest(3)               ",
"/sim_minimips/u_minimips/mem_adr_reg_dest(4)               ",
"/sim_minimips/u_minimips/mem_adr_reg_dest(5)               ",
"/sim_minimips/u_minimips/mem_ecr_reg                       ",
"/sim_minimips/u_minimips/mem_exc_cause(0)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(1)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(2)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(3)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(4)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(5)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(6)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(7)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(8)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(9)                  ",
"/sim_minimips/u_minimips/mem_exc_cause(10)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(11)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(12)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(13)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(14)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(15)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(16)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(17)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(18)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(19)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(20)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(21)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(22)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(23)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(24)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(25)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(26)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(27)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(28)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(29)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(30)                 ",
"/sim_minimips/u_minimips/mem_exc_cause(31)                 ",
"/sim_minimips/u_minimips/mem_level(0)                      ",
"/sim_minimips/u_minimips/mem_level(1)                      ",
"/sim_minimips/u_minimips/mem_it_ok                         ",
"/sim_minimips/u_minimips/write_adr(0)                      ",
"/sim_minimips/u_minimips/write_adr(1)                      ",
"/sim_minimips/u_minimips/write_adr(2)                      ",
"/sim_minimips/u_minimips/write_adr(3)                      ",
"/sim_minimips/u_minimips/write_adr(4)                      ",
"/sim_minimips/u_minimips/write_gpr                         ",
"/sim_minimips/u_minimips/write_scp                         ",
"/sim_minimips/u_minimips/read_adr1(0)                      ",
"/sim_minimips/u_minimips/read_adr1(1)                      ",
"/sim_minimips/u_minimips/read_adr1(2)                      ",
"/sim_minimips/u_minimips/read_adr1(3)                      ",
"/sim_minimips/u_minimips/read_adr1(4)                      ",
"/sim_minimips/u_minimips/read_adr2(0)                      ",
"/sim_minimips/u_minimips/read_adr2(1)                      ",
"/sim_minimips/u_minimips/read_adr2(2)                      ",
"/sim_minimips/u_minimips/read_adr2(3)                      ",
"/sim_minimips/u_minimips/read_adr2(4)                      ",
"/sim_minimips/u_minimips/interrupt                         ",
"/sim_minimips/u_minimips/vecteur_it(0)                     ",
"/sim_minimips/u_minimips/vecteur_it(1)                     ",
"/sim_minimips/u_minimips/vecteur_it(2)                     ",
"/sim_minimips/u_minimips/vecteur_it(3)                     ",
"/sim_minimips/u_minimips/vecteur_it(4)                     ",
"/sim_minimips/u_minimips/vecteur_it(5)                     ",
"/sim_minimips/u_minimips/vecteur_it(6)                     ",
"/sim_minimips/u_minimips/vecteur_it(7)                     ",
"/sim_minimips/u_minimips/vecteur_it(8)                     ",
"/sim_minimips/u_minimips/vecteur_it(9)                     ",
"/sim_minimips/u_minimips/vecteur_it(10)                    ",
"/sim_minimips/u_minimips/vecteur_it(11)                    ",
"/sim_minimips/u_minimips/vecteur_it(12)                    ",
"/sim_minimips/u_minimips/vecteur_it(13)                    ",
"/sim_minimips/u_minimips/vecteur_it(14)                    ",
"/sim_minimips/u_minimips/vecteur_it(15)                    ",
"/sim_minimips/u_minimips/vecteur_it(16)                    ",
"/sim_minimips/u_minimips/vecteur_it(17)                    ",
"/sim_minimips/u_minimips/vecteur_it(18)                    ",
"/sim_minimips/u_minimips/vecteur_it(19)                    ",
"/sim_minimips/u_minimips/vecteur_it(20)                    ",
"/sim_minimips/u_minimips/vecteur_it(21)                    ",
"/sim_minimips/u_minimips/vecteur_it(22)                    ",
"/sim_minimips/u_minimips/vecteur_it(23)                    ",
"/sim_minimips/u_minimips/vecteur_it(24)                    ",
"/sim_minimips/u_minimips/vecteur_it(25)                    ",
"/sim_minimips/u_minimips/vecteur_it(26)                    ",
"/sim_minimips/u_minimips/vecteur_it(27)                    ",
"/sim_minimips/u_minimips/vecteur_it(28)                    ",
"/sim_minimips/u_minimips/vecteur_it(29)                    ",
"/sim_minimips/u_minimips/vecteur_it(30)                    ",
"/sim_minimips/u_minimips/vecteur_it(31)                    ",
"/sim_minimips/u_minimips/pr_bra_bad                        ",
"/sim_minimips/u_minimips/pr_bra_adr(0)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(1)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(2)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(3)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(4)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(5)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(6)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(7)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(8)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(9)                     ",
"/sim_minimips/u_minimips/pr_bra_adr(10)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(11)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(12)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(13)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(14)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(15)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(16)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(17)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(18)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(19)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(20)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(21)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(22)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(23)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(24)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(25)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(26)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(27)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(28)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(29)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(30)                    ",
"/sim_minimips/u_minimips/pr_bra_adr(31)                    ",
"/sim_minimips/u_minimips/pr_clear                          ",
"/sim_minimips/u_minimips/clear                             ",
"/sim_minimips/u_minimips/alea2                             ",
"/sim_minimips/u_minimips/alea3                             ",
"/sim_minimips/u_minimips/u3_di/pre_bra                     ",
"/sim_minimips/u_minimips/u3_di/pre_link                    ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(0)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(1)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(2)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(3)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(4)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(5)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(6)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(7)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(8)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(9)             ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(10)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(11)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(12)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(13)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(14)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(15)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(16)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(17)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(18)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(19)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(20)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(21)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(22)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(23)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(24)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(25)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(26)            ",
"/sim_minimips/u_minimips/u3_di/pre_code_ual(27)            ",
"/sim_minimips/u_minimips/u3_di/pre_offset(0)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(1)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(2)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(3)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(4)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(5)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(6)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(7)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(8)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(9)               ",
"/sim_minimips/u_minimips/u3_di/pre_offset(10)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(11)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(12)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(13)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(14)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(15)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(16)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(17)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(18)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(19)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(20)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(21)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(22)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(23)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(24)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(25)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(26)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(27)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(28)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(29)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(30)              ",
"/sim_minimips/u_minimips/u3_di/pre_offset(31)              ",
"/sim_minimips/u_minimips/u3_di/pre_adr_reg_dest(0)         ",
"/sim_minimips/u_minimips/u3_di/pre_adr_reg_dest(1)         ",
"/sim_minimips/u_minimips/u3_di/pre_adr_reg_dest(2)         ",
"/sim_minimips/u_minimips/u3_di/pre_adr_reg_dest(3)         ",
"/sim_minimips/u_minimips/u3_di/pre_adr_reg_dest(4)         ",
"/sim_minimips/u_minimips/u3_di/pre_adr_reg_dest(5)         ",
"/sim_minimips/u_minimips/u3_di/pre_ecr_reg                 ",
"/sim_minimips/u_minimips/u3_di/pre_mode                    ",
"/sim_minimips/u_minimips/u3_di/pre_op_mem                  ",
"/sim_minimips/u_minimips/u3_di/pre_r_w                     ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(0)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(1)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(2)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(3)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(4)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(5)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(6)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(7)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(8)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(9)            ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(10)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(11)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(12)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(13)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(14)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(15)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(16)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(17)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(18)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(19)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(20)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(21)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(22)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(23)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(24)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(25)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(26)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(27)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(28)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(29)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(30)           ",
"/sim_minimips/u_minimips/u3_di/pre_exc_cause(31)           ",
"/sim_minimips/u_minimips/u3_di/pre_level(0)                ",
"/sim_minimips/u_minimips/u3_di/pre_level(1)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(0)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(1)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(2)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(3)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(4)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(5)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(6)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(7)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(8)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(9)                 ",
"/sim_minimips/u_minimips/u4_ex/base_adr(10)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(11)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(12)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(13)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(14)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(15)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(16)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(17)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(18)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(19)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(20)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(21)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(22)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(23)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(24)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(25)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(26)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(27)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(28)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(29)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(30)                ",
"/sim_minimips/u_minimips/u4_ex/base_adr(31)                ",
"/sim_minimips/u_minimips/u4_ex/pre_ecr_reg                 ",
"/sim_minimips/u_minimips/u4_ex/pre_bra_confirm             ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(0)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(1)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(2)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(3)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(4)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(5)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(6)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(7)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(8)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(9)            ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(10)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(11)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(12)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(13)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(14)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(15)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(16)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(17)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(18)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(19)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(20)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(21)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(22)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(23)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(24)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(25)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(26)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(27)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(28)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(29)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(30)           ",
"/sim_minimips/u_minimips/u4_ex/pre_exc_cause(31)           ",
"/sim_minimips/u_minimips/u4_ex/overflow_ual                ",
"/sim_minimips/u_minimips/u6_renvoi/dep_r1(0)               ",
"/sim_minimips/u_minimips/u6_renvoi/dep_r1(1)               ",
"/sim_minimips/u_minimips/u6_renvoi/dep_r2(0)               ",
"/sim_minimips/u_minimips/u6_renvoi/dep_r2(1)               ",
"/sim_minimips/u_minimips/u6_renvoi/res_reg                 ",
"/sim_minimips/u_minimips/u6_renvoi/res_mem                 ",
"/sim_minimips/u_minimips/u6_renvoi/res_ex                  ",
"/sim_minimips/u_minimips/u6_renvoi/res_di                  ",
"/sim_minimips/u_minimips/u6_renvoi/resolution(0)           ",
"/sim_minimips/u_minimips/u6_renvoi/resolution(1)           ",
"/sim_minimips/u_minimips/u6_renvoi/resolution(2)           ",
"/sim_minimips/u_minimips/u6_renvoi/resolution(3)           ",
"/sim_minimips/u_minimips/u9_bus_ctrl/r_w                   ",
"/sim_minimips/u_minimips/u9_bus_ctrl/req_allowed           "
);
   
  	type list_string2 is array (natural range <> ) of string(1 to 55);
   constant control_signals_gold : list_string2(1 to 911) := 
(
"/sim_minimips/u_gold/u1_pf/suivant(0)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(1)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(2)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(3)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(4)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(5)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(6)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(7)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(8)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(9)                  ",
"/sim_minimips/u_gold/u1_pf/suivant(10)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(11)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(12)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(13)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(14)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(15)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(16)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(17)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(18)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(19)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(20)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(21)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(22)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(23)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(24)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(25)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(26)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(27)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(28)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(29)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(30)                 ",
"/sim_minimips/u_gold/u1_pf/suivant(31)                 ",
"/sim_minimips/u_gold/u1_pf/pc_interne(0)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(1)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(2)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(3)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(4)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(5)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(6)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(7)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(8)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(9)               ",
"/sim_minimips/u_gold/u1_pf/pc_interne(10)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(11)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(12)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(13)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(14)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(15)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(16)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(17)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(18)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(19)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(20)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(21)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(22)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(23)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(24)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(25)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(26)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(27)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(28)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(29)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(30)              ",
"/sim_minimips/u_gold/u1_pf/pc_interne(31)              ",
"/sim_minimips/u_gold/u1_pf/lock                        ",
"/sim_minimips/u_gold/clock                             ",
"/sim_minimips/u_gold/reset                             ",
"/sim_minimips/u_gold/ram_req                           ",
"/sim_minimips/u_gold/ram_adr(0)                        ",
"/sim_minimips/u_gold/ram_adr(1)                        ",
"/sim_minimips/u_gold/ram_adr(2)                        ",
"/sim_minimips/u_gold/ram_adr(3)                        ",
"/sim_minimips/u_gold/ram_adr(4)                        ",
"/sim_minimips/u_gold/ram_adr(5)                        ",
"/sim_minimips/u_gold/ram_adr(6)                        ",
"/sim_minimips/u_gold/ram_adr(7)                        ",
"/sim_minimips/u_gold/ram_adr(8)                        ",
"/sim_minimips/u_gold/ram_adr(9)                        ",
"/sim_minimips/u_gold/ram_adr(10)                       ",
"/sim_minimips/u_gold/ram_adr(11)                       ",
"/sim_minimips/u_gold/ram_adr(12)                       ",
"/sim_minimips/u_gold/ram_adr(13)                       ",
"/sim_minimips/u_gold/ram_adr(14)                       ",
"/sim_minimips/u_gold/ram_adr(15)                       ",
"/sim_minimips/u_gold/ram_adr(16)                       ",
"/sim_minimips/u_gold/ram_adr(17)                       ",
"/sim_minimips/u_gold/ram_adr(18)                       ",
"/sim_minimips/u_gold/ram_adr(19)                       ",
"/sim_minimips/u_gold/ram_adr(20)                       ",
"/sim_minimips/u_gold/ram_adr(21)                       ",
"/sim_minimips/u_gold/ram_adr(22)                       ",
"/sim_minimips/u_gold/ram_adr(23)                       ",
"/sim_minimips/u_gold/ram_adr(24)                       ",
"/sim_minimips/u_gold/ram_adr(25)                       ",
"/sim_minimips/u_gold/ram_adr(26)                       ",
"/sim_minimips/u_gold/ram_adr(27)                       ",
"/sim_minimips/u_gold/ram_adr(28)                       ",
"/sim_minimips/u_gold/ram_adr(29)                       ",
"/sim_minimips/u_gold/ram_adr(30)                       ",
"/sim_minimips/u_gold/ram_adr(31)                       ",
"/sim_minimips/u_gold/ram_r_w                           ",
"/sim_minimips/u_gold/ram_ack                           ",
"/sim_minimips/u_gold/it_mat                            ",
"/sim_minimips/u_gold/stop_all                          ",
"/sim_minimips/u_gold/it_mat_clk                        ",
"/sim_minimips/u_gold/pf_pc(0)                          ",
"/sim_minimips/u_gold/pf_pc(1)                          ",
"/sim_minimips/u_gold/pf_pc(2)                          ",
"/sim_minimips/u_gold/pf_pc(3)                          ",
"/sim_minimips/u_gold/pf_pc(4)                          ",
"/sim_minimips/u_gold/pf_pc(5)                          ",
"/sim_minimips/u_gold/pf_pc(6)                          ",
"/sim_minimips/u_gold/pf_pc(7)                          ",
"/sim_minimips/u_gold/pf_pc(8)                          ",
"/sim_minimips/u_gold/pf_pc(9)                          ",
"/sim_minimips/u_gold/pf_pc(10)                         ",
"/sim_minimips/u_gold/pf_pc(11)                         ",
"/sim_minimips/u_gold/pf_pc(12)                         ",
"/sim_minimips/u_gold/pf_pc(13)                         ",
"/sim_minimips/u_gold/pf_pc(14)                         ",
"/sim_minimips/u_gold/pf_pc(15)                         ",
"/sim_minimips/u_gold/pf_pc(16)                         ",
"/sim_minimips/u_gold/pf_pc(17)                         ",
"/sim_minimips/u_gold/pf_pc(18)                         ",
"/sim_minimips/u_gold/pf_pc(19)                         ",
"/sim_minimips/u_gold/pf_pc(20)                         ",
"/sim_minimips/u_gold/pf_pc(21)                         ",
"/sim_minimips/u_gold/pf_pc(22)                         ",
"/sim_minimips/u_gold/pf_pc(23)                         ",
"/sim_minimips/u_gold/pf_pc(24)                         ",
"/sim_minimips/u_gold/pf_pc(25)                         ",
"/sim_minimips/u_gold/pf_pc(26)                         ",
"/sim_minimips/u_gold/pf_pc(27)                         ",
"/sim_minimips/u_gold/pf_pc(28)                         ",
"/sim_minimips/u_gold/pf_pc(29)                         ",
"/sim_minimips/u_gold/pf_pc(30)                         ",
"/sim_minimips/u_gold/pf_pc(31)                         ",
"/sim_minimips/u_gold/cte_instr(0)                      ",
"/sim_minimips/u_gold/cte_instr(1)                      ",
"/sim_minimips/u_gold/cte_instr(2)                      ",
"/sim_minimips/u_gold/cte_instr(3)                      ",
"/sim_minimips/u_gold/cte_instr(4)                      ",
"/sim_minimips/u_gold/cte_instr(5)                      ",
"/sim_minimips/u_gold/cte_instr(6)                      ",
"/sim_minimips/u_gold/cte_instr(7)                      ",
"/sim_minimips/u_gold/cte_instr(8)                      ",
"/sim_minimips/u_gold/cte_instr(9)                      ",
"/sim_minimips/u_gold/cte_instr(10)                     ",
"/sim_minimips/u_gold/cte_instr(11)                     ",
"/sim_minimips/u_gold/cte_instr(12)                     ",
"/sim_minimips/u_gold/cte_instr(13)                     ",
"/sim_minimips/u_gold/cte_instr(14)                     ",
"/sim_minimips/u_gold/cte_instr(15)                     ",
"/sim_minimips/u_gold/cte_instr(16)                     ",
"/sim_minimips/u_gold/cte_instr(17)                     ",
"/sim_minimips/u_gold/cte_instr(18)                     ",
"/sim_minimips/u_gold/cte_instr(19)                     ",
"/sim_minimips/u_gold/cte_instr(20)                     ",
"/sim_minimips/u_gold/cte_instr(21)                     ",
"/sim_minimips/u_gold/cte_instr(22)                     ",
"/sim_minimips/u_gold/cte_instr(23)                     ",
"/sim_minimips/u_gold/cte_instr(24)                     ",
"/sim_minimips/u_gold/cte_instr(25)                     ",
"/sim_minimips/u_gold/cte_instr(26)                     ",
"/sim_minimips/u_gold/cte_instr(27)                     ",
"/sim_minimips/u_gold/cte_instr(28)                     ",
"/sim_minimips/u_gold/cte_instr(29)                     ",
"/sim_minimips/u_gold/cte_instr(30)                     ",
"/sim_minimips/u_gold/cte_instr(31)                     ",
"/sim_minimips/u_gold/etc_adr(0)                        ",
"/sim_minimips/u_gold/etc_adr(1)                        ",
"/sim_minimips/u_gold/etc_adr(2)                        ",
"/sim_minimips/u_gold/etc_adr(3)                        ",
"/sim_minimips/u_gold/etc_adr(4)                        ",
"/sim_minimips/u_gold/etc_adr(5)                        ",
"/sim_minimips/u_gold/etc_adr(6)                        ",
"/sim_minimips/u_gold/etc_adr(7)                        ",
"/sim_minimips/u_gold/etc_adr(8)                        ",
"/sim_minimips/u_gold/etc_adr(9)                        ",
"/sim_minimips/u_gold/etc_adr(10)                       ",
"/sim_minimips/u_gold/etc_adr(11)                       ",
"/sim_minimips/u_gold/etc_adr(12)                       ",
"/sim_minimips/u_gold/etc_adr(13)                       ",
"/sim_minimips/u_gold/etc_adr(14)                       ",
"/sim_minimips/u_gold/etc_adr(15)                       ",
"/sim_minimips/u_gold/etc_adr(16)                       ",
"/sim_minimips/u_gold/etc_adr(17)                       ",
"/sim_minimips/u_gold/etc_adr(18)                       ",
"/sim_minimips/u_gold/etc_adr(19)                       ",
"/sim_minimips/u_gold/etc_adr(20)                       ",
"/sim_minimips/u_gold/etc_adr(21)                       ",
"/sim_minimips/u_gold/etc_adr(22)                       ",
"/sim_minimips/u_gold/etc_adr(23)                       ",
"/sim_minimips/u_gold/etc_adr(24)                       ",
"/sim_minimips/u_gold/etc_adr(25)                       ",
"/sim_minimips/u_gold/etc_adr(26)                       ",
"/sim_minimips/u_gold/etc_adr(27)                       ",
"/sim_minimips/u_gold/etc_adr(28)                       ",
"/sim_minimips/u_gold/etc_adr(29)                       ",
"/sim_minimips/u_gold/etc_adr(30)                       ",
"/sim_minimips/u_gold/etc_adr(31)                       ",
"/sim_minimips/u_gold/ei_instr(0)                       ",
"/sim_minimips/u_gold/ei_instr(1)                       ",
"/sim_minimips/u_gold/ei_instr(2)                       ",
"/sim_minimips/u_gold/ei_instr(3)                       ",
"/sim_minimips/u_gold/ei_instr(4)                       ",
"/sim_minimips/u_gold/ei_instr(5)                       ",
"/sim_minimips/u_gold/ei_instr(6)                       ",
"/sim_minimips/u_gold/ei_instr(7)                       ",
"/sim_minimips/u_gold/ei_instr(8)                       ",
"/sim_minimips/u_gold/ei_instr(9)                       ",
"/sim_minimips/u_gold/ei_instr(10)                      ",
"/sim_minimips/u_gold/ei_instr(11)                      ",
"/sim_minimips/u_gold/ei_instr(12)                      ",
"/sim_minimips/u_gold/ei_instr(13)                      ",
"/sim_minimips/u_gold/ei_instr(14)                      ",
"/sim_minimips/u_gold/ei_instr(15)                      ",
"/sim_minimips/u_gold/ei_instr(16)                      ",
"/sim_minimips/u_gold/ei_instr(17)                      ",
"/sim_minimips/u_gold/ei_instr(18)                      ",
"/sim_minimips/u_gold/ei_instr(19)                      ",
"/sim_minimips/u_gold/ei_instr(20)                      ",
"/sim_minimips/u_gold/ei_instr(21)                      ",
"/sim_minimips/u_gold/ei_instr(22)                      ",
"/sim_minimips/u_gold/ei_instr(23)                      ",
"/sim_minimips/u_gold/ei_instr(24)                      ",
"/sim_minimips/u_gold/ei_instr(25)                      ",
"/sim_minimips/u_gold/ei_instr(26)                      ",
"/sim_minimips/u_gold/ei_instr(27)                      ",
"/sim_minimips/u_gold/ei_instr(28)                      ",
"/sim_minimips/u_gold/ei_instr(29)                      ",
"/sim_minimips/u_gold/ei_instr(30)                      ",
"/sim_minimips/u_gold/ei_instr(31)                      ",
"/sim_minimips/u_gold/ei_adr(0)                         ",
"/sim_minimips/u_gold/ei_adr(1)                         ",
"/sim_minimips/u_gold/ei_adr(2)                         ",
"/sim_minimips/u_gold/ei_adr(3)                         ",
"/sim_minimips/u_gold/ei_adr(4)                         ",
"/sim_minimips/u_gold/ei_adr(5)                         ",
"/sim_minimips/u_gold/ei_adr(6)                         ",
"/sim_minimips/u_gold/ei_adr(7)                         ",
"/sim_minimips/u_gold/ei_adr(8)                         ",
"/sim_minimips/u_gold/ei_adr(9)                         ",
"/sim_minimips/u_gold/ei_adr(10)                        ",
"/sim_minimips/u_gold/ei_adr(11)                        ",
"/sim_minimips/u_gold/ei_adr(12)                        ",
"/sim_minimips/u_gold/ei_adr(13)                        ",
"/sim_minimips/u_gold/ei_adr(14)                        ",
"/sim_minimips/u_gold/ei_adr(15)                        ",
"/sim_minimips/u_gold/ei_adr(16)                        ",
"/sim_minimips/u_gold/ei_adr(17)                        ",
"/sim_minimips/u_gold/ei_adr(18)                        ",
"/sim_minimips/u_gold/ei_adr(19)                        ",
"/sim_minimips/u_gold/ei_adr(20)                        ",
"/sim_minimips/u_gold/ei_adr(21)                        ",
"/sim_minimips/u_gold/ei_adr(22)                        ",
"/sim_minimips/u_gold/ei_adr(23)                        ",
"/sim_minimips/u_gold/ei_adr(24)                        ",
"/sim_minimips/u_gold/ei_adr(25)                        ",
"/sim_minimips/u_gold/ei_adr(26)                        ",
"/sim_minimips/u_gold/ei_adr(27)                        ",
"/sim_minimips/u_gold/ei_adr(28)                        ",
"/sim_minimips/u_gold/ei_adr(29)                        ",
"/sim_minimips/u_gold/ei_adr(30)                        ",
"/sim_minimips/u_gold/ei_adr(31)                        ",
"/sim_minimips/u_gold/ei_it_ok                          ",
"/sim_minimips/u_gold/adr_reg1(0)                       ",
"/sim_minimips/u_gold/adr_reg1(1)                       ",
"/sim_minimips/u_gold/adr_reg1(2)                       ",
"/sim_minimips/u_gold/adr_reg1(3)                       ",
"/sim_minimips/u_gold/adr_reg1(4)                       ",
"/sim_minimips/u_gold/adr_reg1(5)                       ",
"/sim_minimips/u_gold/adr_reg2(0)                       ",
"/sim_minimips/u_gold/adr_reg2(1)                       ",
"/sim_minimips/u_gold/adr_reg2(2)                       ",
"/sim_minimips/u_gold/adr_reg2(3)                       ",
"/sim_minimips/u_gold/adr_reg2(4)                       ",
"/sim_minimips/u_gold/adr_reg2(5)                       ",
"/sim_minimips/u_gold/use1                              ",
"/sim_minimips/u_gold/use2                              ",
"/sim_minimips/u_gold/alea                              ",
"/sim_minimips/u_gold/di_bra                            ",
"/sim_minimips/u_gold/di_link                           ",
"/sim_minimips/u_gold/di_code_ual(0)                    ",
"/sim_minimips/u_gold/di_code_ual(1)                    ",
"/sim_minimips/u_gold/di_code_ual(2)                    ",
"/sim_minimips/u_gold/di_code_ual(3)                    ",
"/sim_minimips/u_gold/di_code_ual(4)                    ",
"/sim_minimips/u_gold/di_code_ual(5)                    ",
"/sim_minimips/u_gold/di_code_ual(6)                    ",
"/sim_minimips/u_gold/di_code_ual(7)                    ",
"/sim_minimips/u_gold/di_code_ual(8)                    ",
"/sim_minimips/u_gold/di_code_ual(9)                    ",
"/sim_minimips/u_gold/di_code_ual(10)                   ",
"/sim_minimips/u_gold/di_code_ual(11)                   ",
"/sim_minimips/u_gold/di_code_ual(12)                   ",
"/sim_minimips/u_gold/di_code_ual(13)                   ",
"/sim_minimips/u_gold/di_code_ual(14)                   ",
"/sim_minimips/u_gold/di_code_ual(15)                   ",
"/sim_minimips/u_gold/di_code_ual(16)                   ",
"/sim_minimips/u_gold/di_code_ual(17)                   ",
"/sim_minimips/u_gold/di_code_ual(18)                   ",
"/sim_minimips/u_gold/di_code_ual(19)                   ",
"/sim_minimips/u_gold/di_code_ual(20)                   ",
"/sim_minimips/u_gold/di_code_ual(21)                   ",
"/sim_minimips/u_gold/di_code_ual(22)                   ",
"/sim_minimips/u_gold/di_code_ual(23)                   ",
"/sim_minimips/u_gold/di_code_ual(24)                   ",
"/sim_minimips/u_gold/di_code_ual(25)                   ",
"/sim_minimips/u_gold/di_code_ual(26)                   ",
"/sim_minimips/u_gold/di_code_ual(27)                   ",
"/sim_minimips/u_gold/di_offset(0)                      ",
"/sim_minimips/u_gold/di_offset(1)                      ",
"/sim_minimips/u_gold/di_offset(2)                      ",
"/sim_minimips/u_gold/di_offset(3)                      ",
"/sim_minimips/u_gold/di_offset(4)                      ",
"/sim_minimips/u_gold/di_offset(5)                      ",
"/sim_minimips/u_gold/di_offset(6)                      ",
"/sim_minimips/u_gold/di_offset(7)                      ",
"/sim_minimips/u_gold/di_offset(8)                      ",
"/sim_minimips/u_gold/di_offset(9)                      ",
"/sim_minimips/u_gold/di_offset(10)                     ",
"/sim_minimips/u_gold/di_offset(11)                     ",
"/sim_minimips/u_gold/di_offset(12)                     ",
"/sim_minimips/u_gold/di_offset(13)                     ",
"/sim_minimips/u_gold/di_offset(14)                     ",
"/sim_minimips/u_gold/di_offset(15)                     ",
"/sim_minimips/u_gold/di_offset(16)                     ",
"/sim_minimips/u_gold/di_offset(17)                     ",
"/sim_minimips/u_gold/di_offset(18)                     ",
"/sim_minimips/u_gold/di_offset(19)                     ",
"/sim_minimips/u_gold/di_offset(20)                     ",
"/sim_minimips/u_gold/di_offset(21)                     ",
"/sim_minimips/u_gold/di_offset(22)                     ",
"/sim_minimips/u_gold/di_offset(23)                     ",
"/sim_minimips/u_gold/di_offset(24)                     ",
"/sim_minimips/u_gold/di_offset(25)                     ",
"/sim_minimips/u_gold/di_offset(26)                     ",
"/sim_minimips/u_gold/di_offset(27)                     ",
"/sim_minimips/u_gold/di_offset(28)                     ",
"/sim_minimips/u_gold/di_offset(29)                     ",
"/sim_minimips/u_gold/di_offset(30)                     ",
"/sim_minimips/u_gold/di_offset(31)                     ",
"/sim_minimips/u_gold/di_adr_reg_dest(0)                ",
"/sim_minimips/u_gold/di_adr_reg_dest(1)                ",
"/sim_minimips/u_gold/di_adr_reg_dest(2)                ",
"/sim_minimips/u_gold/di_adr_reg_dest(3)                ",
"/sim_minimips/u_gold/di_adr_reg_dest(4)                ",
"/sim_minimips/u_gold/di_adr_reg_dest(5)                ",
"/sim_minimips/u_gold/di_ecr_reg                        ",
"/sim_minimips/u_gold/di_mode                           ",
"/sim_minimips/u_gold/di_op_mem                         ",
"/sim_minimips/u_gold/di_r_w                            ",
"/sim_minimips/u_gold/di_adr(0)                         ",
"/sim_minimips/u_gold/di_adr(1)                         ",
"/sim_minimips/u_gold/di_adr(2)                         ",
"/sim_minimips/u_gold/di_adr(3)                         ",
"/sim_minimips/u_gold/di_adr(4)                         ",
"/sim_minimips/u_gold/di_adr(5)                         ",
"/sim_minimips/u_gold/di_adr(6)                         ",
"/sim_minimips/u_gold/di_adr(7)                         ",
"/sim_minimips/u_gold/di_adr(8)                         ",
"/sim_minimips/u_gold/di_adr(9)                         ",
"/sim_minimips/u_gold/di_adr(10)                        ",
"/sim_minimips/u_gold/di_adr(11)                        ",
"/sim_minimips/u_gold/di_adr(12)                        ",
"/sim_minimips/u_gold/di_adr(13)                        ",
"/sim_minimips/u_gold/di_adr(14)                        ",
"/sim_minimips/u_gold/di_adr(15)                        ",
"/sim_minimips/u_gold/di_adr(16)                        ",
"/sim_minimips/u_gold/di_adr(17)                        ",
"/sim_minimips/u_gold/di_adr(18)                        ",
"/sim_minimips/u_gold/di_adr(19)                        ",
"/sim_minimips/u_gold/di_adr(20)                        ",
"/sim_minimips/u_gold/di_adr(21)                        ",
"/sim_minimips/u_gold/di_adr(22)                        ",
"/sim_minimips/u_gold/di_adr(23)                        ",
"/sim_minimips/u_gold/di_adr(24)                        ",
"/sim_minimips/u_gold/di_adr(25)                        ",
"/sim_minimips/u_gold/di_adr(26)                        ",
"/sim_minimips/u_gold/di_adr(27)                        ",
"/sim_minimips/u_gold/di_adr(28)                        ",
"/sim_minimips/u_gold/di_adr(29)                        ",
"/sim_minimips/u_gold/di_adr(30)                        ",
"/sim_minimips/u_gold/di_adr(31)                        ",
"/sim_minimips/u_gold/di_exc_cause(0)                   ",
"/sim_minimips/u_gold/di_exc_cause(1)                   ",
"/sim_minimips/u_gold/di_exc_cause(2)                   ",
"/sim_minimips/u_gold/di_exc_cause(3)                   ",
"/sim_minimips/u_gold/di_exc_cause(4)                   ",
"/sim_minimips/u_gold/di_exc_cause(5)                   ",
"/sim_minimips/u_gold/di_exc_cause(6)                   ",
"/sim_minimips/u_gold/di_exc_cause(7)                   ",
"/sim_minimips/u_gold/di_exc_cause(8)                   ",
"/sim_minimips/u_gold/di_exc_cause(9)                   ",
"/sim_minimips/u_gold/di_exc_cause(10)                  ",
"/sim_minimips/u_gold/di_exc_cause(11)                  ",
"/sim_minimips/u_gold/di_exc_cause(12)                  ",
"/sim_minimips/u_gold/di_exc_cause(13)                  ",
"/sim_minimips/u_gold/di_exc_cause(14)                  ",
"/sim_minimips/u_gold/di_exc_cause(15)                  ",
"/sim_minimips/u_gold/di_exc_cause(16)                  ",
"/sim_minimips/u_gold/di_exc_cause(17)                  ",
"/sim_minimips/u_gold/di_exc_cause(18)                  ",
"/sim_minimips/u_gold/di_exc_cause(19)                  ",
"/sim_minimips/u_gold/di_exc_cause(20)                  ",
"/sim_minimips/u_gold/di_exc_cause(21)                  ",
"/sim_minimips/u_gold/di_exc_cause(22)                  ",
"/sim_minimips/u_gold/di_exc_cause(23)                  ",
"/sim_minimips/u_gold/di_exc_cause(24)                  ",
"/sim_minimips/u_gold/di_exc_cause(25)                  ",
"/sim_minimips/u_gold/di_exc_cause(26)                  ",
"/sim_minimips/u_gold/di_exc_cause(27)                  ",
"/sim_minimips/u_gold/di_exc_cause(28)                  ",
"/sim_minimips/u_gold/di_exc_cause(29)                  ",
"/sim_minimips/u_gold/di_exc_cause(30)                  ",
"/sim_minimips/u_gold/di_exc_cause(31)                  ",
"/sim_minimips/u_gold/di_level(0)                       ",
"/sim_minimips/u_gold/di_level(1)                       ",
"/sim_minimips/u_gold/di_it_ok                          ",
"/sim_minimips/u_gold/ex_adr(0)                         ",
"/sim_minimips/u_gold/ex_adr(1)                         ",
"/sim_minimips/u_gold/ex_adr(2)                         ",
"/sim_minimips/u_gold/ex_adr(3)                         ",
"/sim_minimips/u_gold/ex_adr(4)                         ",
"/sim_minimips/u_gold/ex_adr(5)                         ",
"/sim_minimips/u_gold/ex_adr(6)                         ",
"/sim_minimips/u_gold/ex_adr(7)                         ",
"/sim_minimips/u_gold/ex_adr(8)                         ",
"/sim_minimips/u_gold/ex_adr(9)                         ",
"/sim_minimips/u_gold/ex_adr(10)                        ",
"/sim_minimips/u_gold/ex_adr(11)                        ",
"/sim_minimips/u_gold/ex_adr(12)                        ",
"/sim_minimips/u_gold/ex_adr(13)                        ",
"/sim_minimips/u_gold/ex_adr(14)                        ",
"/sim_minimips/u_gold/ex_adr(15)                        ",
"/sim_minimips/u_gold/ex_adr(16)                        ",
"/sim_minimips/u_gold/ex_adr(17)                        ",
"/sim_minimips/u_gold/ex_adr(18)                        ",
"/sim_minimips/u_gold/ex_adr(19)                        ",
"/sim_minimips/u_gold/ex_adr(20)                        ",
"/sim_minimips/u_gold/ex_adr(21)                        ",
"/sim_minimips/u_gold/ex_adr(22)                        ",
"/sim_minimips/u_gold/ex_adr(23)                        ",
"/sim_minimips/u_gold/ex_adr(24)                        ",
"/sim_minimips/u_gold/ex_adr(25)                        ",
"/sim_minimips/u_gold/ex_adr(26)                        ",
"/sim_minimips/u_gold/ex_adr(27)                        ",
"/sim_minimips/u_gold/ex_adr(28)                        ",
"/sim_minimips/u_gold/ex_adr(29)                        ",
"/sim_minimips/u_gold/ex_adr(30)                        ",
"/sim_minimips/u_gold/ex_adr(31)                        ",
"/sim_minimips/u_gold/ex_bra_confirm                    ",
"/sim_minimips/u_gold/ex_adresse(0)                     ",
"/sim_minimips/u_gold/ex_adresse(1)                     ",
"/sim_minimips/u_gold/ex_adresse(2)                     ",
"/sim_minimips/u_gold/ex_adresse(3)                     ",
"/sim_minimips/u_gold/ex_adresse(4)                     ",
"/sim_minimips/u_gold/ex_adresse(5)                     ",
"/sim_minimips/u_gold/ex_adresse(6)                     ",
"/sim_minimips/u_gold/ex_adresse(7)                     ",
"/sim_minimips/u_gold/ex_adresse(8)                     ",
"/sim_minimips/u_gold/ex_adresse(9)                     ",
"/sim_minimips/u_gold/ex_adresse(10)                    ",
"/sim_minimips/u_gold/ex_adresse(11)                    ",
"/sim_minimips/u_gold/ex_adresse(12)                    ",
"/sim_minimips/u_gold/ex_adresse(13)                    ",
"/sim_minimips/u_gold/ex_adresse(14)                    ",
"/sim_minimips/u_gold/ex_adresse(15)                    ",
"/sim_minimips/u_gold/ex_adresse(16)                    ",
"/sim_minimips/u_gold/ex_adresse(17)                    ",
"/sim_minimips/u_gold/ex_adresse(18)                    ",
"/sim_minimips/u_gold/ex_adresse(19)                    ",
"/sim_minimips/u_gold/ex_adresse(20)                    ",
"/sim_minimips/u_gold/ex_adresse(21)                    ",
"/sim_minimips/u_gold/ex_adresse(22)                    ",
"/sim_minimips/u_gold/ex_adresse(23)                    ",
"/sim_minimips/u_gold/ex_adresse(24)                    ",
"/sim_minimips/u_gold/ex_adresse(25)                    ",
"/sim_minimips/u_gold/ex_adresse(26)                    ",
"/sim_minimips/u_gold/ex_adresse(27)                    ",
"/sim_minimips/u_gold/ex_adresse(28)                    ",
"/sim_minimips/u_gold/ex_adresse(29)                    ",
"/sim_minimips/u_gold/ex_adresse(30)                    ",
"/sim_minimips/u_gold/ex_adresse(31)                    ",
"/sim_minimips/u_gold/ex_adr_reg_dest(0)                ",
"/sim_minimips/u_gold/ex_adr_reg_dest(1)                ",
"/sim_minimips/u_gold/ex_adr_reg_dest(2)                ",
"/sim_minimips/u_gold/ex_adr_reg_dest(3)                ",
"/sim_minimips/u_gold/ex_adr_reg_dest(4)                ",
"/sim_minimips/u_gold/ex_adr_reg_dest(5)                ",
"/sim_minimips/u_gold/ex_ecr_reg                        ",
"/sim_minimips/u_gold/ex_op_mem                         ",
"/sim_minimips/u_gold/ex_r_w                            ",
"/sim_minimips/u_gold/ex_exc_cause(0)                   ",
"/sim_minimips/u_gold/ex_exc_cause(1)                   ",
"/sim_minimips/u_gold/ex_exc_cause(2)                   ",
"/sim_minimips/u_gold/ex_exc_cause(3)                   ",
"/sim_minimips/u_gold/ex_exc_cause(4)                   ",
"/sim_minimips/u_gold/ex_exc_cause(5)                   ",
"/sim_minimips/u_gold/ex_exc_cause(6)                   ",
"/sim_minimips/u_gold/ex_exc_cause(7)                   ",
"/sim_minimips/u_gold/ex_exc_cause(8)                   ",
"/sim_minimips/u_gold/ex_exc_cause(9)                   ",
"/sim_minimips/u_gold/ex_exc_cause(10)                  ",
"/sim_minimips/u_gold/ex_exc_cause(11)                  ",
"/sim_minimips/u_gold/ex_exc_cause(12)                  ",
"/sim_minimips/u_gold/ex_exc_cause(13)                  ",
"/sim_minimips/u_gold/ex_exc_cause(14)                  ",
"/sim_minimips/u_gold/ex_exc_cause(15)                  ",
"/sim_minimips/u_gold/ex_exc_cause(16)                  ",
"/sim_minimips/u_gold/ex_exc_cause(17)                  ",
"/sim_minimips/u_gold/ex_exc_cause(18)                  ",
"/sim_minimips/u_gold/ex_exc_cause(19)                  ",
"/sim_minimips/u_gold/ex_exc_cause(20)                  ",
"/sim_minimips/u_gold/ex_exc_cause(21)                  ",
"/sim_minimips/u_gold/ex_exc_cause(22)                  ",
"/sim_minimips/u_gold/ex_exc_cause(23)                  ",
"/sim_minimips/u_gold/ex_exc_cause(24)                  ",
"/sim_minimips/u_gold/ex_exc_cause(25)                  ",
"/sim_minimips/u_gold/ex_exc_cause(26)                  ",
"/sim_minimips/u_gold/ex_exc_cause(27)                  ",
"/sim_minimips/u_gold/ex_exc_cause(28)                  ",
"/sim_minimips/u_gold/ex_exc_cause(29)                  ",
"/sim_minimips/u_gold/ex_exc_cause(30)                  ",
"/sim_minimips/u_gold/ex_exc_cause(31)                  ",
"/sim_minimips/u_gold/ex_level(0)                       ",
"/sim_minimips/u_gold/ex_level(1)                       ",
"/sim_minimips/u_gold/ex_it_ok                          ",
"/sim_minimips/u_gold/mtc_adr(0)                        ",
"/sim_minimips/u_gold/mtc_adr(1)                        ",
"/sim_minimips/u_gold/mtc_adr(2)                        ",
"/sim_minimips/u_gold/mtc_adr(3)                        ",
"/sim_minimips/u_gold/mtc_adr(4)                        ",
"/sim_minimips/u_gold/mtc_adr(5)                        ",
"/sim_minimips/u_gold/mtc_adr(6)                        ",
"/sim_minimips/u_gold/mtc_adr(7)                        ",
"/sim_minimips/u_gold/mtc_adr(8)                        ",
"/sim_minimips/u_gold/mtc_adr(9)                        ",
"/sim_minimips/u_gold/mtc_adr(10)                       ",
"/sim_minimips/u_gold/mtc_adr(11)                       ",
"/sim_minimips/u_gold/mtc_adr(12)                       ",
"/sim_minimips/u_gold/mtc_adr(13)                       ",
"/sim_minimips/u_gold/mtc_adr(14)                       ",
"/sim_minimips/u_gold/mtc_adr(15)                       ",
"/sim_minimips/u_gold/mtc_adr(16)                       ",
"/sim_minimips/u_gold/mtc_adr(17)                       ",
"/sim_minimips/u_gold/mtc_adr(18)                       ",
"/sim_minimips/u_gold/mtc_adr(19)                       ",
"/sim_minimips/u_gold/mtc_adr(20)                       ",
"/sim_minimips/u_gold/mtc_adr(21)                       ",
"/sim_minimips/u_gold/mtc_adr(22)                       ",
"/sim_minimips/u_gold/mtc_adr(23)                       ",
"/sim_minimips/u_gold/mtc_adr(24)                       ",
"/sim_minimips/u_gold/mtc_adr(25)                       ",
"/sim_minimips/u_gold/mtc_adr(26)                       ",
"/sim_minimips/u_gold/mtc_adr(27)                       ",
"/sim_minimips/u_gold/mtc_adr(28)                       ",
"/sim_minimips/u_gold/mtc_adr(29)                       ",
"/sim_minimips/u_gold/mtc_adr(30)                       ",
"/sim_minimips/u_gold/mtc_adr(31)                       ",
"/sim_minimips/u_gold/mtc_r_w                           ",
"/sim_minimips/u_gold/mtc_req                           ",
"/sim_minimips/u_gold/mem_adr(0)                        ",
"/sim_minimips/u_gold/mem_adr(1)                        ",
"/sim_minimips/u_gold/mem_adr(2)                        ",
"/sim_minimips/u_gold/mem_adr(3)                        ",
"/sim_minimips/u_gold/mem_adr(4)                        ",
"/sim_minimips/u_gold/mem_adr(5)                        ",
"/sim_minimips/u_gold/mem_adr(6)                        ",
"/sim_minimips/u_gold/mem_adr(7)                        ",
"/sim_minimips/u_gold/mem_adr(8)                        ",
"/sim_minimips/u_gold/mem_adr(9)                        ",
"/sim_minimips/u_gold/mem_adr(10)                       ",
"/sim_minimips/u_gold/mem_adr(11)                       ",
"/sim_minimips/u_gold/mem_adr(12)                       ",
"/sim_minimips/u_gold/mem_adr(13)                       ",
"/sim_minimips/u_gold/mem_adr(14)                       ",
"/sim_minimips/u_gold/mem_adr(15)                       ",
"/sim_minimips/u_gold/mem_adr(16)                       ",
"/sim_minimips/u_gold/mem_adr(17)                       ",
"/sim_minimips/u_gold/mem_adr(18)                       ",
"/sim_minimips/u_gold/mem_adr(19)                       ",
"/sim_minimips/u_gold/mem_adr(20)                       ",
"/sim_minimips/u_gold/mem_adr(21)                       ",
"/sim_minimips/u_gold/mem_adr(22)                       ",
"/sim_minimips/u_gold/mem_adr(23)                       ",
"/sim_minimips/u_gold/mem_adr(24)                       ",
"/sim_minimips/u_gold/mem_adr(25)                       ",
"/sim_minimips/u_gold/mem_adr(26)                       ",
"/sim_minimips/u_gold/mem_adr(27)                       ",
"/sim_minimips/u_gold/mem_adr(28)                       ",
"/sim_minimips/u_gold/mem_adr(29)                       ",
"/sim_minimips/u_gold/mem_adr(30)                       ",
"/sim_minimips/u_gold/mem_adr(31)                       ",
"/sim_minimips/u_gold/mem_adr_reg_dest(0)               ",
"/sim_minimips/u_gold/mem_adr_reg_dest(1)               ",
"/sim_minimips/u_gold/mem_adr_reg_dest(2)               ",
"/sim_minimips/u_gold/mem_adr_reg_dest(3)               ",
"/sim_minimips/u_gold/mem_adr_reg_dest(4)               ",
"/sim_minimips/u_gold/mem_adr_reg_dest(5)               ",
"/sim_minimips/u_gold/mem_ecr_reg                       ",
"/sim_minimips/u_gold/mem_exc_cause(0)                  ",
"/sim_minimips/u_gold/mem_exc_cause(1)                  ",
"/sim_minimips/u_gold/mem_exc_cause(2)                  ",
"/sim_minimips/u_gold/mem_exc_cause(3)                  ",
"/sim_minimips/u_gold/mem_exc_cause(4)                  ",
"/sim_minimips/u_gold/mem_exc_cause(5)                  ",
"/sim_minimips/u_gold/mem_exc_cause(6)                  ",
"/sim_minimips/u_gold/mem_exc_cause(7)                  ",
"/sim_minimips/u_gold/mem_exc_cause(8)                  ",
"/sim_minimips/u_gold/mem_exc_cause(9)                  ",
"/sim_minimips/u_gold/mem_exc_cause(10)                 ",
"/sim_minimips/u_gold/mem_exc_cause(11)                 ",
"/sim_minimips/u_gold/mem_exc_cause(12)                 ",
"/sim_minimips/u_gold/mem_exc_cause(13)                 ",
"/sim_minimips/u_gold/mem_exc_cause(14)                 ",
"/sim_minimips/u_gold/mem_exc_cause(15)                 ",
"/sim_minimips/u_gold/mem_exc_cause(16)                 ",
"/sim_minimips/u_gold/mem_exc_cause(17)                 ",
"/sim_minimips/u_gold/mem_exc_cause(18)                 ",
"/sim_minimips/u_gold/mem_exc_cause(19)                 ",
"/sim_minimips/u_gold/mem_exc_cause(20)                 ",
"/sim_minimips/u_gold/mem_exc_cause(21)                 ",
"/sim_minimips/u_gold/mem_exc_cause(22)                 ",
"/sim_minimips/u_gold/mem_exc_cause(23)                 ",
"/sim_minimips/u_gold/mem_exc_cause(24)                 ",
"/sim_minimips/u_gold/mem_exc_cause(25)                 ",
"/sim_minimips/u_gold/mem_exc_cause(26)                 ",
"/sim_minimips/u_gold/mem_exc_cause(27)                 ",
"/sim_minimips/u_gold/mem_exc_cause(28)                 ",
"/sim_minimips/u_gold/mem_exc_cause(29)                 ",
"/sim_minimips/u_gold/mem_exc_cause(30)                 ",
"/sim_minimips/u_gold/mem_exc_cause(31)                 ",
"/sim_minimips/u_gold/mem_level(0)                      ",
"/sim_minimips/u_gold/mem_level(1)                      ",
"/sim_minimips/u_gold/mem_it_ok                         ",
"/sim_minimips/u_gold/write_adr(0)                      ",
"/sim_minimips/u_gold/write_adr(1)                      ",
"/sim_minimips/u_gold/write_adr(2)                      ",
"/sim_minimips/u_gold/write_adr(3)                      ",
"/sim_minimips/u_gold/write_adr(4)                      ",
"/sim_minimips/u_gold/write_gpr                         ",
"/sim_minimips/u_gold/write_scp                         ",
"/sim_minimips/u_gold/read_adr1(0)                      ",
"/sim_minimips/u_gold/read_adr1(1)                      ",
"/sim_minimips/u_gold/read_adr1(2)                      ",
"/sim_minimips/u_gold/read_adr1(3)                      ",
"/sim_minimips/u_gold/read_adr1(4)                      ",
"/sim_minimips/u_gold/read_adr2(0)                      ",
"/sim_minimips/u_gold/read_adr2(1)                      ",
"/sim_minimips/u_gold/read_adr2(2)                      ",
"/sim_minimips/u_gold/read_adr2(3)                      ",
"/sim_minimips/u_gold/read_adr2(4)                      ",
"/sim_minimips/u_gold/interrupt                         ",
"/sim_minimips/u_gold/vecteur_it(0)                     ",
"/sim_minimips/u_gold/vecteur_it(1)                     ",
"/sim_minimips/u_gold/vecteur_it(2)                     ",
"/sim_minimips/u_gold/vecteur_it(3)                     ",
"/sim_minimips/u_gold/vecteur_it(4)                     ",
"/sim_minimips/u_gold/vecteur_it(5)                     ",
"/sim_minimips/u_gold/vecteur_it(6)                     ",
"/sim_minimips/u_gold/vecteur_it(7)                     ",
"/sim_minimips/u_gold/vecteur_it(8)                     ",
"/sim_minimips/u_gold/vecteur_it(9)                     ",
"/sim_minimips/u_gold/vecteur_it(10)                    ",
"/sim_minimips/u_gold/vecteur_it(11)                    ",
"/sim_minimips/u_gold/vecteur_it(12)                    ",
"/sim_minimips/u_gold/vecteur_it(13)                    ",
"/sim_minimips/u_gold/vecteur_it(14)                    ",
"/sim_minimips/u_gold/vecteur_it(15)                    ",
"/sim_minimips/u_gold/vecteur_it(16)                    ",
"/sim_minimips/u_gold/vecteur_it(17)                    ",
"/sim_minimips/u_gold/vecteur_it(18)                    ",
"/sim_minimips/u_gold/vecteur_it(19)                    ",
"/sim_minimips/u_gold/vecteur_it(20)                    ",
"/sim_minimips/u_gold/vecteur_it(21)                    ",
"/sim_minimips/u_gold/vecteur_it(22)                    ",
"/sim_minimips/u_gold/vecteur_it(23)                    ",
"/sim_minimips/u_gold/vecteur_it(24)                    ",
"/sim_minimips/u_gold/vecteur_it(25)                    ",
"/sim_minimips/u_gold/vecteur_it(26)                    ",
"/sim_minimips/u_gold/vecteur_it(27)                    ",
"/sim_minimips/u_gold/vecteur_it(28)                    ",
"/sim_minimips/u_gold/vecteur_it(29)                    ",
"/sim_minimips/u_gold/vecteur_it(30)                    ",
"/sim_minimips/u_gold/vecteur_it(31)                    ",
"/sim_minimips/u_gold/pr_bra_bad                        ",
"/sim_minimips/u_gold/pr_bra_adr(0)                     ",
"/sim_minimips/u_gold/pr_bra_adr(1)                     ",
"/sim_minimips/u_gold/pr_bra_adr(2)                     ",
"/sim_minimips/u_gold/pr_bra_adr(3)                     ",
"/sim_minimips/u_gold/pr_bra_adr(4)                     ",
"/sim_minimips/u_gold/pr_bra_adr(5)                     ",
"/sim_minimips/u_gold/pr_bra_adr(6)                     ",
"/sim_minimips/u_gold/pr_bra_adr(7)                     ",
"/sim_minimips/u_gold/pr_bra_adr(8)                     ",
"/sim_minimips/u_gold/pr_bra_adr(9)                     ",
"/sim_minimips/u_gold/pr_bra_adr(10)                    ",
"/sim_minimips/u_gold/pr_bra_adr(11)                    ",
"/sim_minimips/u_gold/pr_bra_adr(12)                    ",
"/sim_minimips/u_gold/pr_bra_adr(13)                    ",
"/sim_minimips/u_gold/pr_bra_adr(14)                    ",
"/sim_minimips/u_gold/pr_bra_adr(15)                    ",
"/sim_minimips/u_gold/pr_bra_adr(16)                    ",
"/sim_minimips/u_gold/pr_bra_adr(17)                    ",
"/sim_minimips/u_gold/pr_bra_adr(18)                    ",
"/sim_minimips/u_gold/pr_bra_adr(19)                    ",
"/sim_minimips/u_gold/pr_bra_adr(20)                    ",
"/sim_minimips/u_gold/pr_bra_adr(21)                    ",
"/sim_minimips/u_gold/pr_bra_adr(22)                    ",
"/sim_minimips/u_gold/pr_bra_adr(23)                    ",
"/sim_minimips/u_gold/pr_bra_adr(24)                    ",
"/sim_minimips/u_gold/pr_bra_adr(25)                    ",
"/sim_minimips/u_gold/pr_bra_adr(26)                    ",
"/sim_minimips/u_gold/pr_bra_adr(27)                    ",
"/sim_minimips/u_gold/pr_bra_adr(28)                    ",
"/sim_minimips/u_gold/pr_bra_adr(29)                    ",
"/sim_minimips/u_gold/pr_bra_adr(30)                    ",
"/sim_minimips/u_gold/pr_bra_adr(31)                    ",
"/sim_minimips/u_gold/pr_clear                          ",
"/sim_minimips/u_gold/clear                             ",
"/sim_minimips/u_gold/alea2                             ",
"/sim_minimips/u_gold/alea3                             ",
"/sim_minimips/u_gold/u3_di/pre_bra                     ",
"/sim_minimips/u_gold/u3_di/pre_link                    ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(0)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(1)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(2)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(3)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(4)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(5)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(6)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(7)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(8)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(9)             ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(10)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(11)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(12)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(13)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(14)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(15)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(16)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(17)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(18)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(19)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(20)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(21)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(22)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(23)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(24)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(25)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(26)            ",
"/sim_minimips/u_gold/u3_di/pre_code_ual(27)            ",
"/sim_minimips/u_gold/u3_di/pre_offset(0)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(1)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(2)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(3)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(4)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(5)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(6)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(7)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(8)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(9)               ",
"/sim_minimips/u_gold/u3_di/pre_offset(10)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(11)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(12)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(13)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(14)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(15)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(16)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(17)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(18)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(19)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(20)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(21)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(22)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(23)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(24)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(25)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(26)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(27)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(28)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(29)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(30)              ",
"/sim_minimips/u_gold/u3_di/pre_offset(31)              ",
"/sim_minimips/u_gold/u3_di/pre_adr_reg_dest(0)         ",
"/sim_minimips/u_gold/u3_di/pre_adr_reg_dest(1)         ",
"/sim_minimips/u_gold/u3_di/pre_adr_reg_dest(2)         ",
"/sim_minimips/u_gold/u3_di/pre_adr_reg_dest(3)         ",
"/sim_minimips/u_gold/u3_di/pre_adr_reg_dest(4)         ",
"/sim_minimips/u_gold/u3_di/pre_adr_reg_dest(5)         ",
"/sim_minimips/u_gold/u3_di/pre_ecr_reg                 ",
"/sim_minimips/u_gold/u3_di/pre_mode                    ",
"/sim_minimips/u_gold/u3_di/pre_op_mem                  ",
"/sim_minimips/u_gold/u3_di/pre_r_w                     ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(0)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(1)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(2)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(3)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(4)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(5)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(6)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(7)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(8)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(9)            ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(10)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(11)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(12)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(13)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(14)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(15)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(16)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(17)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(18)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(19)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(20)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(21)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(22)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(23)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(24)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(25)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(26)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(27)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(28)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(29)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(30)           ",
"/sim_minimips/u_gold/u3_di/pre_exc_cause(31)           ",
"/sim_minimips/u_gold/u3_di/pre_level(0)                ",
"/sim_minimips/u_gold/u3_di/pre_level(1)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(0)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(1)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(2)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(3)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(4)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(5)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(6)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(7)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(8)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(9)                 ",
"/sim_minimips/u_gold/u4_ex/base_adr(10)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(11)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(12)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(13)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(14)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(15)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(16)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(17)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(18)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(19)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(20)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(21)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(22)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(23)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(24)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(25)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(26)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(27)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(28)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(29)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(30)                ",
"/sim_minimips/u_gold/u4_ex/base_adr(31)                ",
"/sim_minimips/u_gold/u4_ex/pre_ecr_reg                 ",
"/sim_minimips/u_gold/u4_ex/pre_bra_confirm             ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(0)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(1)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(2)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(3)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(4)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(5)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(6)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(7)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(8)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(9)            ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(10)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(11)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(12)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(13)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(14)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(15)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(16)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(17)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(18)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(19)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(20)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(21)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(22)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(23)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(24)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(25)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(26)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(27)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(28)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(29)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(30)           ",
"/sim_minimips/u_gold/u4_ex/pre_exc_cause(31)           ",
"/sim_minimips/u_gold/u4_ex/overflow_ual                ",
"/sim_minimips/u_gold/u6_renvoi/dep_r1(0)               ",
"/sim_minimips/u_gold/u6_renvoi/dep_r1(1)               ",
"/sim_minimips/u_gold/u6_renvoi/dep_r2(0)               ",
"/sim_minimips/u_gold/u6_renvoi/dep_r2(1)               ",
"/sim_minimips/u_gold/u6_renvoi/res_reg                 ",
"/sim_minimips/u_gold/u6_renvoi/res_mem                 ",
"/sim_minimips/u_gold/u6_renvoi/res_ex                  ",
"/sim_minimips/u_gold/u6_renvoi/res_di                  ",
"/sim_minimips/u_gold/u6_renvoi/resolution(0)           ",
"/sim_minimips/u_gold/u6_renvoi/resolution(1)           ",
"/sim_minimips/u_gold/u6_renvoi/resolution(2)           ",
"/sim_minimips/u_gold/u6_renvoi/resolution(3)           ",
"/sim_minimips/u_gold/u9_bus_ctrl/r_w                   ",
"/sim_minimips/u_gold/u9_bus_ctrl/req_allowed           "
);



  signal reg_uut : std_logic_vector (1 to 992); -- tamanho igual a lista de sinais
  type list_string3 is array (natural range <> ) of string(1 to 50);
  constant reg_signals_uut : list_string3(1 to 992) := 
(
"/sim_minimips/u_minimips/u7_banc/registres(1)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(1)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(2)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(3)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(4)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(5)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(6)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(7)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(8)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(31) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(30) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(29) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(28) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(27) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(26) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(25) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(24) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(23) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(22) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(21) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(20) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(19) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(18) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(17) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(16) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(15) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(14) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(13) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(12) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(11) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(10) ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(9)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(8)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(7)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(6)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(5)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(4)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(3)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(2)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(1)  ",
"/sim_minimips/u_minimips/u7_banc/registres(9)(0)  ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(10)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(10)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(11)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(11)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(12)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(12)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(13)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(13)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(14)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(14)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(15)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(15)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(16)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(16)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(17)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(17)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(18)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(18)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(19)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(19)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(20)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(20)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(21)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(21)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(22)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(22)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(23)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(23)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(24)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(24)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(25)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(25)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(26)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(26)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(27)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(27)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(28)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(28)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(29)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(29)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(30)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(30)(0) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(31)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(30)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(29)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(28)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(27)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(26)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(25)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(24)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(23)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(22)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(21)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(20)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(19)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(18)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(17)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(16)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(15)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(14)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(13)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(12)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(11)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(10)",
"/sim_minimips/u_minimips/u7_banc/registres(31)(9) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(8) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(7) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(6) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(5) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(4) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(3) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(2) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(1) ",
"/sim_minimips/u_minimips/u7_banc/registres(31)(0) "
);

begin

    u_minimips : minimips port map (
        clock => clock,
        reset => reset,
        ram_req => ram_req,
        ram_adr => ram_adr,
        ram_r_w => ram_r_w,
        ram_data => ram_data,
        ram_ack => ram_rdy,
        
        mem_data_out => mem_data_out_in,
        
        it_mat => it_mat
    );

    U_ram : ram port map (
        req => ram_req,
        adr => ram_adr,
        data_inout => ram_data,
        
        --Caco
        mem_data_in => mem_data_out_in,
        
        r_w => ram_r_w,
        ready => ram_rdy,
        reset => reset,
        clock => clock
    );
	
	  --  u_gold : minimips port map (
      --  clock => clock_g,
      --  reset => reset_g,
      --  ram_req => ram_req_g,
      --  ram_adr => ram_adr_g,
      --  ram_r_w => ram_r_w_g,
      --  ram_data => ram_data_g,
      --  ram_ack => ram_rdy_g,
      --  mem_data_out => mem_data_out_in_g,
      --  it_mat => it_mat_g
  --  );

  --  U_ram_gold : ram port map (
  --      req => ram_req_g,
  --      adr => ram_adr_g,
  --      data_inout => ram_data_g,
        
        --Caco
  --      mem_data_in => mem_data_out_in_g,
        
  --      r_w => ram_r_w_g,
  --      ready => ram_rdy_g,
  --      reset => reset_g,
  --      clock => clock_g
  --  );


--   ram_data <= ram_data_temp;
--   ram_data <=  "00000000000000000000000000000000" when end_of_execution='1';

load_signals: process      -- carrega para o sinal forced os sinais da list_signals_1
begin
     for h in 1 to reg_signals_uut'high loop
         init_signal_spy(reg_signals_uut(h),"/sim_minimips/reg_uut(" & integer'image(h)&")",0, 1);
		-- init_signal_spy(reg_signals_gold(h),"/sim_minimips/reg_gold(" & integer'image(h)&")",0, 1);
    end loop;
    wait;
end process;

--load_signals2: process      -- carrega para o sinal forced os sinais da list_signals_1
--begin
--     for h in 1 to control_signals_uut'high loop
--         init_signal_spy(control_signals_uut(h),"/sim_minimips/control_uut(" & integer'image(h)&")",0, 1);
--		 init_signal_spy(control_signals_gold(h),"/sim_minimips/control_gold(" & integer'image(h)&")",0, 1);
--    end loop;
--    wait;
--end process;



process
begin
clock <= '0';
clock_g <= '0';
wait for 21 ns;
clock <= '1';
clock_g <= '1';
wait for 21 ns;
end process;


--    ram_data <= (others => 'L');

   -- END OF EXECUTION
   process (ram_adr, clock)
    begin 
       if (ram_adr = "00000000000000000000000111101100") then
             debug1 <= '1';
       else
             debug1 <= '0';
       end if;
    end process;
   
   
    process (ram_adr)
    begin 
        --if (ram_r_w = '1') then
--       if (ram_adr = "00000000000000000000001000001100") then -- teste2
--       if (ram_adr = "00000000000000000000001001110100") then -- teste4
  --if (ram_adr = "00000000000000000000001010001100") then -- bubble10
  --if (ram_adr = "00000000000000000000001010001100") then -- bubble20
									   
     --  if (ram_adr = "00000000000000000000001011101100") then -- select10
--       if (ram_adr = "00000000000000000000001011101100") then -- select3
--       if (ram_adr = "00000000000000000000001111111100") then -- quick10
--       if (ram_adr = "00000000000000000000010101000100") then -- imdct

--       if (ram_adr = "00000000000000000000011111011000") then -- stringsearch
--         if (ram_adr = "00000000000000000000001010111000") then -- select_teste
                                      
 --if (ram_adr = "00000000000000000000001001000000") then -- testeFuncao
-- if (ram_adr = "00000000000000000000010001011000") then ---quick100_mips2.coe
if (ram_adr = "00000000000000000000001110110000") then ---quick_mips.coe
									 
            end_of_execution <= '1';
         end if;
    end process;

    process (ram_adr_g, clock_g)
    begin 
       if (ram_adr_g = "00000000000000000000000111101100") then
             debug1_g <= '1';
       else
             debug1_g <= '0';
       end if;
    end process;
	
    process (ram_adr_g)
    begin 
        --if (ram_r_w = '1') then
--       if (ram_adr = "00000000000000000000001000001100") then -- teste2
--       if (ram_adr = "00000000000000000000001001110100") then -- teste4
  --if (ram_adr = "00000000000000000000001010001100") then -- bubble10
  --if (ram_adr = "00000000000000000000001010001100") then -- bubble20
									   
     --  if (ram_adr = "00000000000000000000001011101100") then -- select10
--       if (ram_adr = "00000000000000000000001011101100") then -- select3
--       if (ram_adr = "00000000000000000000001111111100") then -- quick10
--       if (ram_adr = "00000000000000000000010101000100") then -- imdct

--       if (ram_adr = "00000000000000000000011111011000") then -- stringsearch
--         if (ram_adr = "00000000000000000000001010111000") then -- select_teste
                                      
 --if (ram_adr = "00000000000000000000001001000000") then -- testeFuncao
-- if (ram_adr = "00000000000000000000010001011000") then ---quick100_mips2.coe
if (ram_adr = "00000000000000000000001110110000") then ---quick_mips.coe
									 
            end_of_execution_g <= '1';
         end if;
    end process;

    process 
	variable txt1 : line;
	variable txt2 : line;
	variable txt3 : line;
	file fsim1 : text open append_mode is "results.txt";
	file fsim3 : text open append_mode is "counters.txt";
	file fsim2 : text open append_mode is "relatorio.txt";
	variable countFaults: integer:=0;		--number of every faults inserted
	variable failure: integer:=0;		--number of every faults inserted
	variable noeffect : integer:=0;
	variable falhaocorreu : integer := 0;
	variable teste: integer := 0;
	
   begin
  -- while true loop
      reset <= '1';
	  reset_g <= '1';
      wait for 70 ns;
      reset <= '0';
	  reset_g <= '0';
	  countFaults:= countFaults + 1;
	  falhaocorreu := 0;
     wait for 1236263 ns;  --1st 
		
				write (txt1, string'("Falha "));      --place output signals
				write(txt1, countFaults);
				
				write (txt2, string'("Falha "));      --place output signals
				write(txt2, countFaults);
				
				write (txt3, string'("Falha "));      --place output signals
				write(txt3, countFaults);
				
				writeline(fsim2, txt2);
				
				write (txt1, string'(" time: "));		
				write(txt1, string'(integer'image(integer(to_real(now)))));
				write (txt1, string'("ns"));
				
				write (txt3, string'(" time: "));		
				write(txt3, string'(integer'image(integer(to_real(now)))));
				write (txt3, string'("ns"));
				
				if (reg_uut = "00000000010011111111000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000010100000000000000000000000000000101") then
				falhaocorreu := 0;
				
				write (txt2, string'(" Resultado 1 Correto - "));      --place output signals
				--write(txt2, teste);
				
				else
				
				write (txt2, string'(" Resultado 1 Errado - "));      --place output signals
				write(txt2, str(reg_uut));
				falhaocorreu := falhaocorreu +1;
		
				end if;
				
	
				
	wait for 2646 ns;  --2nd 2646  1238979
	
	         if (reg_uut = "00000000010011111111000000000000000000000000000000000000000001010000000000000000000000000000010100000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100") then
	
				write (txt2, string'("Resultado 2 Correto - "));      --place output signals
				--write(txt2, teste);
				
				else
				
				write (txt2, string'("Resultado 2 Errado - "));      --place output signals
				write(txt2, str(reg_uut));
				falhaocorreu := falhaocorreu +1;
				end if;
				
	wait for 2646 ns;  --3rd 1241625
	
	         if (reg_uut = "00000000010011111111000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000010100000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000010101000000000000000000000000000101010000000000000000000000000001010100000000000000000000000000010101000000000000000000000000000101010000000000000000000000000001010100000000000000000000000000101010000000000000000000000000001010100000000000000000000000000010101000000000000000000000000000101010000000000000000000000000001010100000000000000000000000000010101000000000000000000000000000111111000000000000000000000000001111110000000000000000000000000011111100000000000000000000000000111111") then
	
				write (txt2, string'("Resultado 3 Correto - "));      --place output signals
				--write(txt2, teste);
				
				else
				
				write (txt2, string'("Resultado 3 Errado - "));      --place output signals
				write(txt2, str(reg_uut));
				falhaocorreu := falhaocorreu +1;
				end if;
				
   wait for 2058 ns;  --4th  1243683
	
	         if (reg_uut(1 to 768) = "000000000100111111110000000000000000000000000000000000000011111100000000000000000000000000111111000000000000000000000000010101000000000000000000000000000101010000000000000000000000000001010100000000000000000000000000010101000000000000000000000000000101010000000000000000000000000001010100000000000000000000000000011010010000000000000000000000000110100100000000000000000000000001101001000000000000000000000000011010010000000000000000000000000110100100000000000000000000000001101001000000000000000000000000011111100000000000000000000000000111111000000000000000000000000001111110000000000000000000000000011111100000000000000000000000000111111000000000000000000000000001111110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110") then
	
				write (txt2, string'("Resultado 4 Correto"));      --place output signals
				
				else
				
				write (txt2, string'("Resultado 4 Errado"));      --place output signals
				write(txt2, str(reg_uut(1 to 768)));
				falhaocorreu := falhaocorreu +1;
				end if;
				
    writeline(fsim2, txt2);
    
    if (falhaocorreu = 0) then
        write (txt1, string'(" - - Resultado Final Correto")); 
        noeffect := noeffect +1; 
    else
            write (txt1, string'(" - - Resultado Final Errado"));  
            failure := failure + 1;
   end if;
         
     writeline(fsim1, txt1);
	 write (txt3, string'(" NoEffect: "));  
     write(txt3, noeffect);
	 
	  write (txt3, string'(" failure: "));  
     write(txt3, failure);
	 
	 writeline(fsim3, txt3);
   --  end loop;
    wait;
    end process;
	

--process (control_uut, control_gold)
--	variable txt : line;
--	variable txt2 : line;
--	file fsim : text open write_mode is "resultscontrole.txt";
--	file fsim2 : text open write_mode is "reportcontrole.txt";
--begin
	
--	if (clock = '1' and clock'event) then
--	if (control_uut /= control_gold) then
	
--	for i in 1 to control_signals_uut'high loop
--	if (control_uut(i) /= control_gold(i)) then
--		write (txt2, control_signals_gold(i));
--		write (txt2, string'(" "));      --colocar tbm os valores dos sinais
		
 --   end if;
--	end loop;
		
--		write (txt, string'("time: "));		
--		write(txt, string'(integer'image(integer(to_real(now)))));
--		write (txt, string'("ns"));
--		write (txt, string'(" uut: "));	
--		write(txt, str(control_uut));
--		write (txt, string'(" gold: "));	
--		write(txt, str(control_gold));
--		writeline(fsim, txt);
--		writeline(fsim2, txt2);
 --    end if;
--	 end if;
--end process;
	

--    process (ram_adr, ram_r_w, ram_data)
--    begin -- Emulation of an I/O controller
--        ram_data <= (others => 'Z');

--        case ram_adr is
--            when X"00001000" => -- declenche une lecture avec interruption
--                                it_mat <= '1' after 1000 ns;
--                                ram_rdy <= '1' after 5 ns;
--            when X"00001001" => -- fournit la donnee et lache l'it
--                                it_mat <= '0';
--                                ram_data <= X"FFFFFFFF";
--                                ram_rdy <= '1' after 5 ns;
--            when others      => ram_rdy <= 'L';
--        end case;
--    end process;

end bench;




// IVB checksum: 2148765629

`define UFRGS_MINIMIPS_KIT_VERSION "09.20-FIXME"
`define UFRGS_MINIMIPS_KIT_DATE "2009-09-??-FIXME"

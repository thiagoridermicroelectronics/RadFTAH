// IVB checksum: 3210198659
/*-----------------------------------------------------------------
File name     : UFRGS_miniMIPS_types.sv
Developers    : traugusto
Created       : Sun Mar  8 01:06:00 2015
Description   :
Notes         :
-------------------------------------------------------------------
Copyright 2015 (c) Universidade Federal do Rio Grande do Sul
-----------------------------------------------------------------*/

//------------------------------------------------------------------------------
//
// UFRGS_miniMIPS type definitions: enums, parameters, etc
//
//------------------------------------------------------------------------------

typedef enum { NOP,
               READ,
               WRITE
             } UFRGS_miniMIPS_read_write_enum;

